 module _synth_100 (
    input i1,
    input [25 : 0] i2,
    input i3,
    input [31 : 0] i4,
    output [35 : 0] o1
 );
 ADDSUB inst_1(.i1({1'b0, i4[31:0], 3'b000}),
              .i2({9'b000000000, i2[25:0], i3}),
              .i3(i1),
              .o1(o1[35:0]));
 endmodule

 module ADDSUB (
    input [35 : 0] i1,
    input [35 : 0] i2,
    input i3,
    output [35 : 0] o1
 );
 QQ inst_1(.i1(i3),
          .i2(i1[35:0]),
          .i3(i2[35:0]),
          .o1(o1[35:0]));
 endmodule

 module QQ (
    input i1,
    input [35 : 0] i2,
    input [35 : 0] i3,
    output [35 : 0] o1
 );
 wire m188;
 wire m1;
 wire m2;
 wire m3;
 wire m15;
 wire m27;
 wire m32;
 wire m33;
 wire m34;
 wire m35;
 wire m36;
 wire m37;
 wire m38;
 wire m39;
 wire m40;
 wire m41;
 wire m42;
 wire m43;
 wire m44;
 wire m45;
 wire m46;
 wire m4;
 wire m5;
 wire m6;
 wire m7;
 wire m8;
 wire m9;
 wire m10;
 wire m11;
 wire m12;
 wire m13;
 wire m14;
 wire m16;
 wire m17;
 wire m18;
 wire m19;
 wire m20;
 wire m21;
 wire m22;
 wire m23;
 wire m24;
 wire m25;
 wire m26;
 wire m28;
 wire m29;
 wire m30;
 wire m31;
 wire m47;
 wire m48;
 wire m49;
 wire m50;
 wire m51;
 wire m52;
 wire m53;
 wire m85;
 wire m86;
 wire m87;
 wire m88;
 wire m89;
 wire m90;
 wire m91;
 wire m92;
 wire m93;
 wire m94;
 wire m95;
 wire m96;
 wire m97;
 wire m98;
 wire m99;
 wire m100;
 wire m101;
 wire m102;
 wire m103;
 wire m104;
 wire m105;
 wire m106;
 wire m107;
 wire m108;
 wire m109;
 wire m110;
 wire m111;
 wire m112;
 wire m113;
 wire m114;
 wire m115;
 wire m116;
 wire m117;
 wire m118;
 wire m119;
 wire m120;
 wire m54;
 wire m55;
 wire m56;
 wire m57;
 wire m58;
 wire m59;
 wire m60;
 wire m61;
 wire m62;
 wire m63;
 wire m64;
 wire m65;
 wire m66;
 wire m67;
 wire m68;
 wire m69;
 wire m70;
 wire m71;
 wire m72;
 wire m73;
 wire m74;
 wire m75;
 wire m76;
 wire m77;
 wire m78;
 wire m79;
 wire m80;
 wire m81;
 wire m82;
 wire m83;
 wire m84;
 wire m121;
 wire m122;
 wire m123;
 wire m124;
 wire m125;
 wire m142;
 wire m143;
 wire m144;
 wire m145;
 wire m146;
 wire m147;
 wire m148;
 wire m149;
 wire m150;
 wire m151;
 wire m152;
 wire m153;
 wire m154;
 wire m155;
 wire m156;
 wire m157;
 wire m158;
 wire m159;
 wire m160;
 wire m161;
 wire m162;
 wire m163;
 wire m164;
 wire m165;
 wire m166;
 wire m167;
 wire m168;
 wire m169;
 wire m170;
 wire m171;
 wire m172;
 wire m173;
 wire m174;
 wire m175;
 wire m176;
 wire m177;
 wire m178;
 wire m179;
 wire m180;
 wire m181;
 wire m182;
 wire m126;
 wire m127;
 wire m128;
 wire m129;
 wire m130;
 wire m131;
 wire m132;
 wire m133;
 wire m134;
 wire m135;
 wire m136;
 wire m137;
 wire m138;
 wire m139;
 wire m140;
 wire m141;
 wire m183;
 wire m184;
 wire m185;
 wire m186;
 wire m187;
 m_15 inst_1(.i1(i2[0]),
            .i2(m3),
            .i3(i3[0]),
            .o1(m188));
 m_9 inst_2(.i1(m188),
           .i2(m126),
           .i3(m1),
           .o1(m57));
 m_10 inst_3(.i1(i3[35]),
            .i2(i2[35]),
            .o1(m2));
 m_11 inst_4(.i1(i1),
            .o1(m3));
 m_4 inst_5(.i1(i1),
           .i2(m2),
           .o1(m47));
 m_4 inst_6(.i1(i1),
           .i2(i3[34]),
           .o1(m15));
 m_4 inst_7(.i1(i1),
           .i2(i3[2]),
           .o1(m4));
 m_3 inst_8(.i1(i2[2]),
           .i2(m4),
           .o1(m181));
 m_4 inst_9(.i1(i1),
           .i2(i3[3]),
           .o1(m5));
 m_12 inst_10(.i1(i2[3]),
             .i2(m5),
             .o1(m179));
 m_4 inst_11(.i1(i1),
            .i2(i3[4]),
            .o1(m6));
 m_3 inst_12(.i1(i2[4]),
            .i2(m6),
            .o1(m176));
 m_4 inst_13(.i1(i1),
            .i2(i3[5]),
            .o1(m7));
 m_12 inst_14(.i1(i2[5]),
             .i2(m7),
             .o1(m174));
 m_4 inst_15(.i1(i1),
            .i2(i3[6]),
            .o1(m8));
 m_3 inst_16(.i1(i2[6]),
            .i2(m8),
            .o1(m171));
 m_4 inst_17(.i1(i1),
            .i2(i3[7]),
            .o1(m9));
 m_12 inst_18(.i1(i2[7]),
             .i2(m9),
             .o1(m169));
 m_4 inst_19(.i1(i1),
            .i2(i3[8]),
            .o1(m10));
 m_3 inst_20(.i1(i2[8]),
            .i2(m10),
            .o1(m166));
 m_4 inst_21(.i1(i1),
            .i2(i3[9]),
            .o1(m11));
 m_12 inst_22(.i1(i2[9]),
             .i2(m11),
             .o1(m164));
 m_4 inst_23(.i1(i1),
            .i2(i3[10]),
            .o1(m12));
 m_12 inst_24(.i1(i2[10]),
             .i2(m12),
             .o1(m113));
 m_3 inst_25(.i1(i2[10]),
            .i2(m12),
            .o1(m13));
 m_4 inst_26(.i1(i1),
            .i2(i3[11]),
            .o1(m14));
 m_12 inst_27(.i1(i2[11]),
             .i2(m14),
             .o1(m160));
 m_6 inst_28(.i1(i2[34]),
            .i2(m15),
            .o1(m61));
 m_3 inst_29(.i1(i2[34]),
            .i2(m15),
            .o1(m65));
 m_4 inst_30(.i1(i1),
            .i2(i3[33]),
            .o1(m27));
 m_4 inst_31(.i1(i1),
            .i2(i3[12]),
            .o1(m16));
 m_3 inst_32(.i1(i2[12]),
            .i2(m16),
            .o1(m109));
 m_4 inst_33(.i1(i1),
            .i2(i3[13]),
            .o1(m17));
 m_4 inst_34(.i1(i1),
            .i2(i3[14]),
            .o1(m18));
 m_3 inst_35(.i1(i2[14]),
            .i2(m18),
            .o1(m100));
 m_4 inst_36(.i1(i1),
            .i2(i3[15]),
            .o1(m19));
 m_4 inst_37(.i1(i1),
            .i2(i3[16]),
            .o1(m20));
 m_12 inst_38(.i1(i2[16]),
             .i2(m20),
             .o1(m92));
 m_10 inst_39(.i1(i2[16]),
             .i2(m20),
             .o1(m156));
 m_4 inst_40(.i1(i1),
            .i2(i3[17]),
            .o1(m21));
 m_12 inst_41(.i1(i2[17]),
             .i2(m21),
             .o1(m90));
 m_3 inst_42(.i1(i2[17]),
            .i2(m21),
            .o1(m22));
 m_4 inst_43(.i1(i1),
            .i2(i3[18]),
            .o1(m23));
 m_6 inst_44(.i1(i2[18]),
            .i2(m23),
            .o1(m148));
 m_4 inst_45(.i1(i1),
            .i2(i3[19]),
            .o1(m24));
 m_6 inst_46(.i1(i2[19]),
            .i2(m24),
            .o1(m151));
 m_13 inst_47(.i1(i2[19]),
             .i2(m24),
             .o1(m145));
 m_4 inst_48(.i1(i1),
            .i2(i3[20]),
            .o1(m25));
 m_6 inst_49(.i1(i2[20]),
            .i2(m25),
            .o1(m86));
 m_4 inst_50(.i1(i1),
            .i2(i3[21]),
            .o1(m26));
 m_6 inst_51(.i1(i2[21]),
            .i2(m26),
            .o1(m88));
 m_13 inst_52(.i1(i2[21]),
             .i2(m26),
             .o1(m186));
 m_13 inst_53(.i1(i2[33]),
             .i2(m27),
             .o1(m67));
 m_4 inst_54(.i1(i1),
            .i2(i3[32]),
            .o1(m32));
 m_4 inst_55(.i1(i1),
            .i2(i3[22]),
            .o1(m28));
 m_6 inst_56(.i1(i2[22]),
            .i2(m28),
            .o1(m122));
 m_4 inst_57(.i1(i1),
            .i2(i3[23]),
            .o1(m29));
 m_6 inst_58(.i1(i2[23]),
            .i2(m29),
            .o1(m124));
 m_13 inst_59(.i1(i2[23]),
             .i2(m29),
             .o1(m125));
 m_4 inst_60(.i1(i1),
            .i2(i3[24]),
            .o1(m30));
 m_12 inst_61(.i1(i2[24]),
             .i2(m30),
             .o1(m31));
 m_4 inst_62(.i1(i2[24]),
            .i2(m30),
            .o1(m138));
 m_6 inst_63(.i1(i2[32]),
            .i2(m32),
            .o1(m33));
 m_13 inst_64(.i1(i2[32]),
             .i2(m32),
             .o1(m34));
 m_4 inst_65(.i1(i1),
            .i2(i3[31]),
            .o1(m35));
 m_13 inst_66(.i1(i2[31]),
             .i2(m35),
             .o1(m131));
 m_4 inst_67(.i1(i1),
            .i2(i3[30]),
            .o1(m36));
 m_6 inst_68(.i1(i2[30]),
            .i2(m36),
            .o1(m74));
 m_13 inst_69(.i1(i2[30]),
             .i2(m36),
             .o1(m75));
 m_4 inst_70(.i1(i1),
            .i2(i3[29]),
            .o1(m37));
 m_6 inst_71(.i1(i2[29]),
            .i2(m37),
            .o1(m38));
 m_13 inst_72(.i1(i2[29]),
             .i2(m37),
             .o1(m39));
 m_8 inst_73(.i1(m53),
            .i2(m133),
            .i3(m39),
            .o1(m77));
 m_4 inst_74(.i1(i1),
            .i2(i3[27]),
            .o1(m40));
 m_12 inst_75(.i1(i2[27]),
             .i2(m40),
             .o1(m41));
 m_3 inst_76(.i1(i2[27]),
            .i2(m40),
            .o1(m42));
 m_4 inst_77(.i1(i1),
            .i2(i3[26]),
            .o1(m43));
 m_12 inst_78(.i1(i2[26]),
             .i2(m43),
             .o1(m44));
 m_6 inst_79(.i1(m44),
            .i2(m41),
            .o1(m45));
 m_4 inst_80(.i1(i2[26]),
            .i2(m43),
            .o1(m136));
 m_4 inst_81(.i1(i1),
            .i2(i3[1]),
            .o1(m46));
 m_12 inst_82(.i1(i2[1]),
             .i2(m46),
             .o1(m1));
 m_4 inst_83(.i1(i2[1]),
            .i2(m46),
            .o1(m126));
 m_4 inst_84(.i1(i3[25]),
            .i2(i1),
            .o1(m48));
 m_12 inst_85(.i1(i2[25]),
             .i2(m48),
             .o1(m49));
 m_12 inst_86(.i1(m31),
             .i2(m49),
             .o1(m51));
 m_3 inst_87(.i1(i2[25]),
            .i2(m48),
            .o1(m50));
 m_9 inst_88(.i1(m139),
            .i2(m51),
            .i3(m50),
            .o1(m137));
 m_10 inst_89(.i1(i1),
             .i2(i3[28]),
             .o1(m52));
 m_3 inst_90(.i1(m79),
            .i2(m52),
            .o1(m53));
 m_4 inst_91(.i1(m121),
            .i2(m123),
            .o1(o1[23]));
 m_4 inst_92(.i1(m85),
            .i2(m87),
            .o1(o1[21]));
 m_4 inst_93(.i1(m54),
            .i2(m55),
            .o1(o1[4]));
 m_12 inst_94(.i1(m56),
             .i2(m176),
             .o1(m55));
 m_12 inst_95(.i1(i2[4]),
             .i2(m6),
             .o1(m56));
 m_4 inst_96(.i1(m57),
            .i2(m58),
            .o1(o1[2]));
 m_12 inst_97(.i1(m59),
             .i2(m181),
             .o1(m58));
 m_12 inst_98(.i1(i2[2]),
             .i2(m4),
             .o1(m59));
 m_4 inst_99(.i1(m60),
            .i2(m47),
            .o1(o1[35]));
 m_8 inst_100(.i1(m62),
             .i2(m65),
             .i3(m61),
             .o1(m60));
 m_4 inst_101(.i1(m62),
             .i2(m63),
             .o1(o1[34]));
 m_12 inst_102(.i1(m64),
              .i2(m65),
              .o1(m63));
 m_12 inst_103(.i1(i2[34]),
              .i2(m15),
              .o1(m64));
 m_4 inst_104(.i1(m66),
             .i2(m69),
             .o1(o1[33]));
 m_9 inst_105(.i1(m66),
             .i2(m67),
             .i3(m68),
             .o1(m62));
 m_12 inst_106(.i1(i2[33]),
              .i2(m27),
              .o1(m68));
 m_10 inst_107(.i1(i2[33]),
              .i2(m27),
              .o1(m69));
 m_4 inst_108(.i1(m70),
             .i2(m72),
             .o1(o1[31]));
 m_9 inst_109(.i1(m75),
             .i2(m76),
             .i3(m71),
             .o1(m70));
 m_12 inst_110(.i1(i2[30]),
              .i2(m36),
              .o1(m71));
 m_4 inst_111(.i1(i2[31]),
             .i2(m35),
             .o1(m72));
 m_4 inst_112(.i1(m73),
             .i2(m76),
             .o1(o1[30]));
 m_13 inst_113(.i1(m74),
              .i2(m75),
              .o1(m73));
 m_9 inst_114(.i1(m38),
             .i2(m77),
             .i3(m73),
             .o1(m129));
 m_13 inst_115(.i1(m38),
              .i2(m77),
              .o1(m76));
 m_4 inst_116(.i1(m78),
             .i2(m80),
             .o1(o1[29]));
 m_9 inst_117(.i1(m79),
             .i2(m52),
             .i3(m133),
             .o1(m78));
 m_11 inst_118(.i1(i2[28]),
              .o1(m79));
 m_3 inst_119(.i1(m38),
             .i2(m39),
             .o1(m80));
 m_4 inst_120(.i1(m81),
             .i2(m82),
             .o1(o1[27]));
 m_9 inst_121(.i1(m136),
             .i2(m137),
             .i3(m44),
             .o1(m81));
 m_12 inst_122(.i1(m41),
              .i2(m42),
              .o1(m82));
 m_4 inst_123(.i1(m83),
             .i2(m84),
             .o1(o1[25]));
 m_9 inst_124(.i1(m138),
             .i2(m140),
             .i3(m31),
             .o1(m83));
 m_12 inst_125(.i1(m49),
              .i2(m50),
              .o1(m84));
 m_3 inst_126(.i1(m86),
             .i2(m143),
             .o1(m85));
 m_3 inst_127(.i1(m88),
             .i2(m186),
             .o1(m87));
 m_4 inst_128(.i1(m89),
             .i2(m91),
             .o1(o1[17]));
 m_12 inst_129(.i1(m22),
              .i2(m90),
              .o1(m89));
 m_12 inst_130(.i1(m92),
              .i2(m93),
              .o1(m91));
 m_12 inst_131(.i1(m92),
              .i2(m90),
              .o1(m157));
 m_4 inst_132(.i1(m94),
             .i2(m97),
             .o1(o1[15]));
 m_9 inst_133(.i1(m95),
             .i2(m94),
             .i3(m96),
             .o1(m158));
 m_13 inst_134(.i1(i2[15]),
              .i2(m19),
              .o1(m95));
 m_12 inst_135(.i1(i2[15]),
              .i2(m19),
              .o1(m96));
 m_10 inst_136(.i1(i2[15]),
              .i2(m19),
              .o1(m97));
 m_4 inst_137(.i1(m98),
             .i2(m101),
             .o1(o1[14]));
 m_12 inst_138(.i1(m99),
              .i2(m100),
              .o1(m98));
 m_12 inst_139(.i1(i2[14]),
              .i2(m18),
              .o1(m99));
 m_8 inst_140(.i1(m100),
             .i2(m101),
             .i3(m102),
             .o1(m94));
 m_6 inst_141(.i1(i2[14]),
             .i2(m18),
             .o1(m102));
 m_4 inst_142(.i1(m103),
             .i2(m106),
             .o1(o1[13]));
 m_9 inst_143(.i1(m104),
             .i2(m103),
             .i3(m105),
             .o1(m101));
 m_13 inst_144(.i1(i2[13]),
              .i2(m17),
              .o1(m104));
 m_12 inst_145(.i1(i2[13]),
              .i2(m17),
              .o1(m105));
 m_10 inst_146(.i1(i2[13]),
              .i2(m17),
              .o1(m106));
 m_4 inst_147(.i1(m107),
             .i2(m110),
             .o1(o1[12]));
 m_12 inst_148(.i1(m108),
              .i2(m109),
              .o1(m107));
 m_12 inst_149(.i1(i2[12]),
              .i2(m16),
              .o1(m108));
 m_8 inst_150(.i1(m109),
             .i2(m110),
             .i3(m111),
             .o1(m103));
 m_6 inst_151(.i1(i2[12]),
             .i2(m16),
             .o1(m111));
 m_4 inst_152(.i1(m112),
             .i2(m114),
             .o1(o1[10]));
 m_12 inst_153(.i1(m113),
              .i2(m13),
              .o1(m112));
 m_4 inst_154(.i1(m115),
             .i2(m116),
             .o1(o1[8]));
 m_12 inst_155(.i1(m117),
              .i2(m166),
              .o1(m116));
 m_12 inst_156(.i1(i2[8]),
              .i2(m10),
              .o1(m117));
 m_4 inst_157(.i1(m118),
             .i2(m120),
             .o1(o1[6]));
 m_12 inst_158(.i1(m119),
              .i2(m171),
              .o1(m118));
 m_12 inst_159(.i1(i2[6]),
              .i2(m8),
              .o1(m119));
 m_3 inst_160(.i1(m122),
             .i2(m184),
             .o1(m121));
 m_3 inst_161(.i1(m124),
             .i2(m125),
             .o1(m123));
 m inst_162(.i1(m124),
           .i2(m122),
           .i3(m184),
           .o1(m141));
 m_10 inst_163(.i1(m183),
              .i2(m185),
              .o1(o1[22]));
 m_10 inst_164(.i1(m142),
              .i2(m144),
              .o1(o1[20]));
 m_10 inst_165(.i1(m188),
              .i2(m126),
              .o1(o1[1]));
 m_10 inst_166(.i1(i3[0]),
              .i2(i2[0]),
              .o1(o1[0]));
 m_10 inst_167(.i1(m127),
              .i2(m128),
              .o1(o1[32]));
 m_8 inst_168(.i1(m127),
             .i2(m128),
             .i3(m33),
             .o1(m66));
 m_13 inst_169(.i1(m33),
              .i2(m34),
              .o1(m127));
 m_8 inst_170(.i1(m129),
             .i2(m130),
             .i3(m131),
             .o1(m128));
 m_8 inst_171(.i1(i2[31]),
             .i2(m35),
             .i3(m74),
             .o1(m130));
 m_10 inst_172(.i1(m132),
              .i2(m134),
              .o1(o1[28]));
 m_14 inst_173(.i1(m42),
              .i2(m132),
              .i3(m135),
              .o1(m133));
 m_4 inst_174(.i1(i2[28]),
             .i2(m52),
             .o1(m132));
 m_6 inst_175(.i1(m42),
             .i2(m135),
             .o1(m134));
 m_9 inst_176(.i1(m136),
             .i2(m137),
             .i3(m45),
             .o1(m135));
 m_10 inst_177(.i1(m136),
              .i2(m137),
              .o1(o1[26]));
 m_10 inst_178(.i1(m138),
              .i2(m140),
              .o1(o1[24]));
 m inst_179(.i1(m138),
           .i2(m125),
           .i3(m141),
           .o1(m139));
 m_3 inst_180(.i1(m125),
             .i2(m141),
             .o1(m140));
 m inst_181(.i1(m142),
           .i2(m145),
           .i3(m146),
           .o1(m143));
 m_4 inst_182(.i1(i2[20]),
             .i2(m25),
             .o1(m142));
 m_3 inst_183(.i1(m145),
             .i2(m146),
             .o1(m144));
 m_10 inst_184(.i1(m147),
              .i2(m150),
              .o1(o1[19]));
 m_3 inst_185(.i1(m148),
             .i2(m149),
             .o1(m147));
 m inst_186(.i1(m151),
           .i2(m148),
           .i3(m149),
           .o1(m146));
 m_13 inst_187(.i1(m151),
              .i2(m145),
              .o1(m150));
 m_10 inst_188(.i1(m152),
              .i2(m153),
              .o1(o1[18]));
 m inst_189(.i1(m152),
           .i2(m154),
           .i3(m155),
           .o1(m149));
 m_4 inst_190(.i1(i2[18]),
             .i2(m23),
             .o1(m152));
 m_3 inst_191(.i1(m154),
             .i2(m155),
             .o1(m153));
 m_11 inst_192(.i1(m22),
              .o1(m154));
 m_10 inst_193(.i1(m156),
              .i2(m158),
              .o1(o1[16]));
 m_8 inst_194(.i1(m156),
             .i2(m158),
             .i3(m157),
             .o1(m155));
 m_12 inst_195(.i1(m156),
              .i2(m158),
              .o1(m93));
 m_10 inst_196(.i1(m159),
              .i2(m161),
              .o1(o1[11]));
 m_9 inst_197(.i1(m159),
             .i2(m161),
             .i3(m160),
             .o1(m110));
 m_4 inst_198(.i1(i2[11]),
             .i2(m14),
             .o1(m159));
 m_8 inst_199(.i1(m13),
             .i2(m114),
             .i3(m162),
             .o1(m161));
 m_11 inst_200(.i1(m113),
              .o1(m162));
 m_10 inst_201(.i1(m163),
              .i2(m165),
              .o1(o1[9]));
 m_9 inst_202(.i1(m163),
             .i2(m165),
             .i3(m164),
             .o1(m114));
 m_4 inst_203(.i1(i2[9]),
             .i2(m11),
             .o1(m163));
 m_8 inst_204(.i1(m115),
             .i2(m166),
             .i3(m167),
             .o1(m165));
 m_6 inst_205(.i1(i2[8]),
             .i2(m10),
             .o1(m167));
 m_10 inst_206(.i1(m168),
              .i2(m170),
              .o1(o1[7]));
 m_9 inst_207(.i1(m168),
             .i2(m170),
             .i3(m169),
             .o1(m115));
 m_4 inst_208(.i1(i2[7]),
             .i2(m9),
             .o1(m168));
 m_8 inst_209(.i1(m171),
             .i2(m120),
             .i3(m172),
             .o1(m170));
 m_6 inst_210(.i1(i2[6]),
             .i2(m8),
             .o1(m172));
 m_10 inst_211(.i1(m173),
              .i2(m175),
              .o1(o1[5]));
 m_9 inst_212(.i1(m173),
             .i2(m175),
             .i3(m174),
             .o1(m120));
 m_4 inst_213(.i1(i2[5]),
             .i2(m7),
             .o1(m173));
 m_8 inst_214(.i1(m54),
             .i2(m176),
             .i3(m177),
             .o1(m175));
 m_6 inst_215(.i1(i2[4]),
             .i2(m6),
             .o1(m177));
 m_10 inst_216(.i1(m178),
              .i2(m180),
              .o1(o1[3]));
 m_9 inst_217(.i1(m178),
             .i2(m180),
             .i3(m179),
             .o1(m54));
 m_4 inst_218(.i1(i2[3]),
             .i2(m5),
             .o1(m178));
 m_8 inst_219(.i1(m57),
             .i2(m181),
             .i3(m182),
             .o1(m180));
 m_6 inst_220(.i1(i2[2]),
             .i2(m4),
             .o1(m182));
 m inst_221(.i1(m183),
           .i2(m186),
           .i3(m187),
           .o1(m184));
 m_4 inst_222(.i1(i2[22]),
             .i2(m28),
             .o1(m183));
 m_3 inst_223(.i1(m186),
             .i2(m187),
             .o1(m185));
 m inst_224(.i1(m88),
           .i2(m86),
           .i3(m143),
           .o1(m187));
 endmodule

 module m_15 (
    input i1,
    input i2,
    input i3,
    output o1
 );
 wire m1;
 m_16 inst_1(.i1(i3),
            .i2(i1),
            .i3(i2),
            .o1(m1));
 m_2 inst_2(.i1(m1),
           .o1(o1));
 endmodule

 module m_16 (
    input i1,
    input i2,
    input i3,
    output o1
 );
 assign o1 = i1 ? i2 : i3;
 endmodule

 module m_14 (
    input i1,
    input i2,
    input i3,
    output o1
 );
 wire m1;
 wire m2;
 m_2 inst_1(.i1(m2),
           .o1(o1));
 m_7 inst_2(.i1(m1),
           .i2(i3),
           .o1(m2));
 m_7 inst_3(.i1(i1),
           .i2(i2),
           .o1(m1));
 endmodule

 module m_13 (
    input i1,
    input i2,
    output o1
 );
 wire m1;
 m_2 inst_1(.i1(m1),
           .o1(o1));
 m_1 inst_2(.i1(i1),
           .i2(i2),
           .o1(m1));
 endmodule

 module m_12 (
    input i1,
    input i2,
    output o1
 );
 wire m1;
 m_2 inst_1(.i1(m1),
           .o1(o1));
 m_7 inst_2(.i1(i1),
           .i2(i2),
           .o1(m1));
 endmodule

 module m_11 (
    input i1,
    output o1
 );
 m_2 inst_1(.i1(i1),
           .o1(o1));
 endmodule

 module m_10 (
    input i1,
    input i2,
    output o1
 );
 m_5 inst_1(.i1(i1),
           .i2(i2),
           .o1(o1));
 endmodule

 module m_9 (
    input i1,
    input i2,
    input i3,
    output o1
 );
 wire m1;
 wire m2;
 m_2 inst_1(.i1(m1),
           .o1(o1));
 m_7 inst_2(.i1(m2),
           .i2(i3),
           .o1(m1));
 m_1 inst_3(.i1(i1),
           .i2(i2),
           .o1(m2));
 endmodule

 module m_8 (
    input i1,
    input i2,
    input i3,
    output o1
 );
 wire m1;
 wire m2;
 m_2 inst_1(.i1(m1),
           .o1(o1));
 m_1 inst_2(.i1(m2),
           .i2(i3),
           .o1(m1));
 m_7 inst_3(.i1(i1),
           .i2(i2),
           .o1(m2));
 endmodule

 module m_6 (
    input i1,
    input i2,
    output o1
 );
 m_7 inst_1(.i1(i1),
           .i2(i2),
           .o1(o1));
 endmodule

 module m_7 (
    input i1,
    input i2,
    output o1
 );
 assign o1 = i1 & i2;
 endmodule

 module m_4 (
    input i1,
    input i2,
    output o1
 );
 wire m1;
 m_2 inst_1(.i1(m1),
           .o1(o1));
 m_5 inst_2(.i1(i1),
           .i2(i2),
           .o1(m1));
 endmodule

 module m_5 (
    input i1,
    input i2,
    output o1
 );
 assign o1 = ~(i1) & i2 | i1 & ~(i2);
 endmodule

 module m_3 (
    input i1,
    input i2,
    output o1
 );
 m_1 inst_1(.i1(i1),
           .i2(i2),
           .o1(o1));
 endmodule

 module m (
    input i1,
    input i2,
    input i3,
    output o1
 );
 wire m1;
 wire m2;
 m_2 inst_1(.i1(m2),
           .o1(o1));
 m_1 inst_2(.i1(m1),
           .i2(i3),
           .o1(m2));
 m_1 inst_3(.i1(i1),
           .i2(i2),
           .o1(m1));
 endmodule

 module m_2 (
    input i1,
    output o1
 );
 assign o1 = ~(i1);
 endmodule

 module m_1 (
    input i1,
    input i2,
    output o1
 );
 assign o1 = i1 | i2;
 endmodule

