 module _synth_106 (
    input [1 : 0] i1,
    input [1 : 0] i2,
    input [3 : 0] i3,
    input [31 : 0] i4,
    input [31 : 0] i5,
    input [33 : 0] i6,
    input [31 : 0] i7,
    input [35 : 0] i8,
    input [1 : 0] i9,
    input [33 : 0] i10,
    input [33 : 0] i11,
    input [1 : 0] i12,
    input i13,
    input i14,
    input [8 : 0] i15,
    input i16,
    input i17,
    input [33 : 0] i18,
    input i19,
    output [36 : 0] o1,
    output [1 : 0] o2,
    output o3,
    output [19 : 0] o4,
    output [33 : 0] o5,
    output [31 : 0] o6,
    output [34 : 0] o7,
    output o8,
    output o9,
    output [8 : 0] o10,
    output o11,
    output o12,
    output o13,
    output o14,
    output [10 : 0] o15,
    output o16,
    output o17,
    output [30 : 0] o18,
    output o19,
    output o20,
    output [24 : 0] o21,
    output [24 : 0] o22
 );
 wire m5;
 wire [1 : 0] m1;
 wire [1 : 0] m2;
 wire m3;
 wire m4;
 Comb inst_1(.i1(i1[1:0]),
            .i2(i2[1:0]),
            .i3(i3[3:0]),
            .i4(i4[31:0]),
            .i5(i5[31:0]),
            .i6(i6[33:0]),
            .i7(i7[31:0]),
            .i8({i8[35:34], m5, i8[33:0]}),
            .i9(i9[1:0]),
            .i10({i10[33:0], m1[1:0]}),
            .i11({i11[33:0], m2[1:0]}),
            .i12(i12[1:0]),
            .i13(i13),
            .i14(i14),
            .i15({m3, i15[8:0]}),
            .i16(i16),
            .i17(i17),
            .i18({i18[33:0], m4}),
            .i19(i19),
            .o1(o1[36:0]),
            .o2(o3),
            .o3(o4[19:0]),
            .o4(o5[33:0]),
            .o5(o6[31:0]),
            .o6(o7[34:0]),
            .o7(o8),
            .o8(o9),
            .o9(o10[8:0]),
            .o10(o11),
            .o11(o12),
            .o12(o13),
            .o13(o14),
            .o14({o15[10:0], o2[1:0]}),
            .o15(o16),
            .o16(o17),
            .o17(o18[30:0]),
            .o18(o19),
            .o19(o20),
            .o20(o21[24:0]),
            .o21(o22[24:0]));
 m_1 inst_2(.i1(1'b0),
           .o1(m5));
 m_1 inst_3(.i1(1'b0),
           .o1(m3));
 m_1 inst_4(.i1(o17),
           .o1(m4));
 m inst_5(.i1(2'b00),
         .o1(m1[1:0]));
 m inst_6(.i1(2'b00),
         .o1(m2[1:0]));
 endmodule

 module Comb (
    input [1 : 0] i1,
    input [1 : 0] i2,
    input [3 : 0] i3,
    input [31 : 0] i4,
    input [31 : 0] i5,
    input [33 : 0] i6,
    input [31 : 0] i7,
    input [36 : 0] i8,
    input [1 : 0] i9,
    input [35 : 0] i10,
    input [35 : 0] i11,
    input [1 : 0] i12,
    input i13,
    input i14,
    input [9 : 0] i15,
    input i16,
    input i17,
    input [34 : 0] i18,
    input i19,
    output [36 : 0] o1,
    output o2,
    output [19 : 0] o3,
    output [33 : 0] o4,
    output [31 : 0] o5,
    output [34 : 0] o6,
    output o7,
    output o8,
    output [8 : 0] o9,
    output o10,
    output o11,
    output o12,
    output o13,
    output [12 : 0] o14,
    output o15,
    output o16,
    output [30 : 0] o17,
    output o18,
    output o19,
    output [24 : 0] o20,
    output [24 : 0] o21
 );
 wire m182;
 wire m183;
 wire m184;
 wire m185;
 wire m186;
 wire m187;
 wire m188;
 wire m189;
 wire m190;
 wire m191;
 wire m192;
 wire m193;
 wire m194;
 wire m195;
 wire m196;
 wire m197;
 wire m198;
 wire m199;
 wire m200;
 wire m201;
 wire m202;
 wire m203;
 wire m204;
 wire m205;
 wire m206;
 wire m207;
 wire m208;
 wire m209;
 wire m210;
 wire m211;
 wire m212;
 wire m213;
 wire m214;
 wire m215;
 wire m216;
 wire m217;
 wire m218;
 wire m219;
 wire m220;
 wire m221;
 wire m222;
 wire m223;
 wire m224;
 wire m225;
 wire m226;
 wire m227;
 wire m228;
 wire m229;
 wire m230;
 wire m231;
 wire m1461;
 wire m1;
 wire m2;
 wire m3;
 wire m4;
 wire m5;
 wire m6;
 wire m7;
 wire m8;
 wire m9;
 wire m10;
 wire m11;
 wire m12;
 wire m13;
 wire m14;
 wire m15;
 wire m16;
 wire m17;
 wire m18;
 wire m19;
 wire m20;
 wire m21;
 wire m22;
 wire m23;
 wire m24;
 wire m25;
 wire m26;
 wire m27;
 wire m28;
 wire m29;
 wire m30;
 wire m31;
 wire m32;
 wire m33;
 wire m34;
 wire m35;
 wire m36;
 wire m37;
 wire m38;
 wire m39;
 wire m40;
 wire m41;
 wire m42;
 wire m43;
 wire m44;
 wire m45;
 wire m46;
 wire m47;
 wire m48;
 wire m49;
 wire m50;
 wire m51;
 wire m52;
 wire m53;
 wire m54;
 wire m55;
 wire m56;
 wire m57;
 wire m58;
 wire m59;
 wire m60;
 wire m61;
 wire m62;
 wire m63;
 wire m64;
 wire m65;
 wire m66;
 wire m67;
 wire m68;
 wire m69;
 wire m70;
 wire m71;
 wire m72;
 wire m73;
 wire m74;
 wire m75;
 wire m76;
 wire m77;
 wire m78;
 wire m79;
 wire m80;
 wire m81;
 wire m82;
 wire m83;
 wire m84;
 wire m85;
 wire m86;
 wire m87;
 wire m88;
 wire m89;
 wire m90;
 wire m91;
 wire m92;
 wire m93;
 wire m94;
 wire m95;
 wire m96;
 wire m97;
 wire m98;
 wire m99;
 wire m100;
 wire m101;
 wire m102;
 wire m103;
 wire m104;
 wire m105;
 wire m106;
 wire m107;
 wire m108;
 wire m109;
 wire m110;
 wire m111;
 wire m112;
 wire m113;
 wire m114;
 wire m115;
 wire m116;
 wire m117;
 wire m118;
 wire m119;
 wire m120;
 wire m121;
 wire m122;
 wire m123;
 wire m124;
 wire m125;
 wire m126;
 wire m127;
 wire m128;
 wire m129;
 wire m130;
 wire m131;
 wire m132;
 wire m133;
 wire m134;
 wire m135;
 wire m136;
 wire m137;
 wire m138;
 wire m139;
 wire m140;
 wire m141;
 wire m142;
 wire m143;
 wire m144;
 wire m145;
 wire m146;
 wire m147;
 wire m148;
 wire m149;
 wire m150;
 wire m151;
 wire m152;
 wire m153;
 wire m154;
 wire m155;
 wire m156;
 wire m157;
 wire m158;
 wire m159;
 wire m160;
 wire m161;
 wire m162;
 wire m163;
 wire m164;
 wire m165;
 wire m166;
 wire m167;
 wire m168;
 wire m169;
 wire m170;
 wire m171;
 wire m172;
 wire m173;
 wire m174;
 wire m175;
 wire m176;
 wire m177;
 wire m178;
 wire m179;
 wire m180;
 wire m181;
 wire m1202;
 wire m1203;
 wire m1204;
 wire m1205;
 wire m1206;
 wire m1207;
 wire m1208;
 wire m1209;
 wire m1210;
 wire m1211;
 wire m1212;
 wire m1213;
 wire m1214;
 wire m1215;
 wire m1216;
 wire m1217;
 wire m1218;
 wire m1219;
 wire m1220;
 wire m1221;
 wire m1222;
 wire m1223;
 wire m1224;
 wire m1225;
 wire m1226;
 wire m1227;
 wire m1228;
 wire m1229;
 wire m1230;
 wire m1231;
 wire m1232;
 wire m1233;
 wire m1234;
 wire m1235;
 wire m1236;
 wire m1237;
 wire m1238;
 wire m1239;
 wire m1240;
 wire m1241;
 wire m1242;
 wire m1243;
 wire m1244;
 wire m1245;
 wire m1246;
 wire m1247;
 wire m1248;
 wire m1249;
 wire m1250;
 wire m1251;
 wire m1252;
 wire m1253;
 wire m1254;
 wire m1255;
 wire m1256;
 wire m1257;
 wire m1258;
 wire m1259;
 wire m1260;
 wire m1261;
 wire m1262;
 wire m1263;
 wire m1264;
 wire m1265;
 wire m1266;
 wire m1267;
 wire m1268;
 wire m1269;
 wire m1270;
 wire m1271;
 wire m1272;
 wire m1273;
 wire m1274;
 wire m1275;
 wire m1276;
 wire m1277;
 wire m1278;
 wire m1279;
 wire m1280;
 wire m1281;
 wire m1282;
 wire m1283;
 wire m1284;
 wire m1285;
 wire m1286;
 wire m1287;
 wire m1288;
 wire m1289;
 wire m1290;
 wire m1291;
 wire m1292;
 wire m1293;
 wire m1294;
 wire m1295;
 wire m1296;
 wire m1297;
 wire m1298;
 wire m1299;
 wire m1300;
 wire m1301;
 wire m1302;
 wire m1303;
 wire m1304;
 wire m1305;
 wire m1306;
 wire m1307;
 wire m1308;
 wire m1309;
 wire m1310;
 wire m1311;
 wire m1312;
 wire m1313;
 wire m1314;
 wire m1315;
 wire m1316;
 wire m1317;
 wire m1318;
 wire m1319;
 wire m1320;
 wire m1321;
 wire m1322;
 wire m1323;
 wire m1324;
 wire m1325;
 wire m1326;
 wire m1357;
 wire m1358;
 wire m1359;
 wire m1369;
 wire m1370;
 wire m1371;
 wire m1372;
 wire m1373;
 wire m1374;
 wire m1375;
 wire m1376;
 wire m1377;
 wire m1378;
 wire m1379;
 wire m1380;
 wire m1381;
 wire m1382;
 wire m1383;
 wire m1384;
 wire m1385;
 wire m1386;
 wire m1387;
 wire m1388;
 wire m1389;
 wire m1390;
 wire m1391;
 wire m1392;
 wire m1327;
 wire m1328;
 wire m1329;
 wire m1330;
 wire m1331;
 wire m1332;
 wire m1333;
 wire m1334;
 wire m1335;
 wire m1336;
 wire m1337;
 wire m1338;
 wire m1339;
 wire m1340;
 wire m1341;
 wire m1342;
 wire m1343;
 wire m1344;
 wire m1345;
 wire m1346;
 wire m1347;
 wire m1348;
 wire m1349;
 wire m1350;
 wire m1351;
 wire m1352;
 wire m1353;
 wire m1354;
 wire m1355;
 wire m1356;
 wire m1360;
 wire m1361;
 wire m1362;
 wire m1363;
 wire m1364;
 wire m1365;
 wire m1366;
 wire m1367;
 wire m1368;
 wire m1393;
 wire m1394;
 wire m1395;
 wire m1396;
 wire m1397;
 wire m1398;
 wire m1399;
 wire m1400;
 wire m1401;
 wire m1402;
 wire m1403;
 wire m1404;
 wire m1405;
 wire m1406;
 wire m1407;
 wire m1408;
 wire m1409;
 wire m1410;
 wire m1411;
 wire m1412;
 wire m1413;
 wire m1414;
 wire m1415;
 wire m1416;
 wire m1417;
 wire m1418;
 wire m1419;
 wire m1420;
 wire m1421;
 wire m1422;
 wire m1423;
 wire m1424;
 wire m1435;
 wire m1439;
 wire m1440;
 wire m1441;
 wire m1442;
 wire m1443;
 wire m1444;
 wire m1445;
 wire m1446;
 wire m1425;
 wire m1426;
 wire m1427;
 wire m1428;
 wire m1429;
 wire m1430;
 wire m1431;
 wire m1432;
 wire m1433;
 wire m1434;
 wire m1436;
 wire m1437;
 wire m1438;
 wire m1447;
 wire m1448;
 wire m1449;
 wire m1450;
 wire m1451;
 wire m1452;
 wire m1453;
 wire m1454;
 wire m1455;
 wire m1456;
 wire m1457;
 wire m1458;
 wire m1459;
 wire m1460;
 wire m232;
 wire m233;
 wire m234;
 wire m235;
 wire m236;
 wire m237;
 wire m238;
 wire m239;
 wire m240;
 wire m241;
 wire m242;
 wire m243;
 wire m244;
 wire m245;
 wire m246;
 wire m247;
 wire m248;
 wire m249;
 wire m250;
 wire m251;
 wire m252;
 wire m253;
 wire m254;
 wire m255;
 wire m256;
 wire m257;
 wire m258;
 wire m259;
 wire m260;
 wire m261;
 wire m262;
 wire m263;
 wire m264;
 wire m265;
 wire m266;
 wire m267;
 wire m268;
 wire m269;
 wire m270;
 wire m271;
 wire m272;
 wire m273;
 wire m274;
 wire m275;
 wire m276;
 wire m277;
 wire m278;
 wire m279;
 wire m280;
 wire m281;
 wire m282;
 wire m283;
 wire m284;
 wire m285;
 wire m286;
 wire m287;
 wire m288;
 wire m289;
 wire m290;
 wire m291;
 wire m292;
 wire m293;
 wire m294;
 wire m295;
 wire m296;
 wire m297;
 wire m298;
 wire m299;
 wire m300;
 wire m301;
 wire m302;
 wire m303;
 wire m304;
 wire m305;
 wire m306;
 wire m307;
 wire m308;
 wire m309;
 wire m310;
 wire m311;
 wire m312;
 wire m313;
 wire m314;
 wire m315;
 wire m316;
 wire m317;
 wire m318;
 wire m319;
 wire m320;
 wire m321;
 wire m322;
 wire m323;
 wire m324;
 wire m325;
 wire m326;
 wire m327;
 wire m328;
 wire m329;
 wire m330;
 wire m331;
 wire m332;
 wire m333;
 wire m334;
 wire m335;
 wire m336;
 wire m337;
 wire m338;
 wire m339;
 wire m340;
 wire m341;
 wire m342;
 wire m343;
 wire m344;
 wire m345;
 wire m346;
 wire m347;
 wire m348;
 wire m349;
 wire m350;
 wire m351;
 wire m352;
 wire m353;
 wire m354;
 wire m355;
 wire m356;
 wire m357;
 wire m358;
 wire m359;
 wire m360;
 wire m361;
 wire m362;
 wire m363;
 wire m364;
 wire m365;
 wire m366;
 wire m367;
 wire m368;
 wire m369;
 wire m370;
 wire m371;
 wire m372;
 wire m373;
 wire m374;
 wire m375;
 wire m376;
 wire m377;
 wire m378;
 wire m379;
 wire m380;
 wire m381;
 wire m382;
 wire m383;
 wire m384;
 wire m385;
 wire m386;
 wire m387;
 wire m388;
 wire m389;
 wire m390;
 wire m391;
 wire m392;
 wire m393;
 wire m394;
 wire m395;
 wire m396;
 wire m397;
 wire m398;
 wire m399;
 wire m400;
 wire m401;
 wire m402;
 wire m403;
 wire m404;
 wire m405;
 wire m406;
 wire m407;
 wire m408;
 wire m409;
 wire m410;
 wire m411;
 wire m412;
 wire m413;
 wire m414;
 wire m415;
 wire m416;
 wire m417;
 wire m418;
 wire m419;
 wire m420;
 wire m421;
 wire m422;
 wire m423;
 wire m424;
 wire m425;
 wire m426;
 wire m427;
 wire m428;
 wire m429;
 wire m430;
 wire m431;
 wire m432;
 wire m433;
 wire m434;
 wire m435;
 wire m436;
 wire m437;
 wire m438;
 wire m439;
 wire m440;
 wire m441;
 wire m442;
 wire m443;
 wire m444;
 wire m445;
 wire m446;
 wire m447;
 wire m448;
 wire m449;
 wire m450;
 wire m451;
 wire m452;
 wire m453;
 wire m454;
 wire m455;
 wire m456;
 wire m457;
 wire m458;
 wire m459;
 wire m460;
 wire m461;
 wire m462;
 wire m463;
 wire m464;
 wire m465;
 wire m466;
 wire m467;
 wire m468;
 wire m469;
 wire m470;
 wire m471;
 wire m472;
 wire m473;
 wire m474;
 wire m475;
 wire m476;
 wire m477;
 wire m478;
 wire m479;
 wire m480;
 wire m481;
 wire m482;
 wire m483;
 wire m484;
 wire m485;
 wire m486;
 wire m487;
 wire m488;
 wire m489;
 wire m490;
 wire m491;
 wire m492;
 wire m493;
 wire m494;
 wire m495;
 wire m496;
 wire m497;
 wire m498;
 wire m499;
 wire m500;
 wire m501;
 wire m502;
 wire m503;
 wire m504;
 wire m505;
 wire m506;
 wire m507;
 wire m508;
 wire m509;
 wire m510;
 wire m511;
 wire m512;
 wire m513;
 wire m514;
 wire m515;
 wire m516;
 wire m517;
 wire m518;
 wire m519;
 wire m520;
 wire m521;
 wire m522;
 wire m523;
 wire m524;
 wire m525;
 wire m526;
 wire m527;
 wire m528;
 wire m529;
 wire m530;
 wire m531;
 wire m532;
 wire m533;
 wire m534;
 wire m535;
 wire m536;
 wire m537;
 wire m538;
 wire m539;
 wire m540;
 wire m541;
 wire m542;
 wire m543;
 wire m544;
 wire m545;
 wire m546;
 wire m547;
 wire m548;
 wire m549;
 wire m550;
 wire m551;
 wire m552;
 wire m553;
 wire m554;
 wire m555;
 wire m556;
 wire m557;
 wire m558;
 wire m559;
 wire m560;
 wire m561;
 wire m562;
 wire m563;
 wire m564;
 wire m565;
 wire m566;
 wire m567;
 wire m568;
 wire m569;
 wire m570;
 wire m571;
 wire m572;
 wire m573;
 wire m574;
 wire m575;
 wire m576;
 wire m577;
 wire m578;
 wire m579;
 wire m580;
 wire m581;
 wire m582;
 wire m583;
 wire m584;
 wire m585;
 wire m586;
 wire m587;
 wire m588;
 wire m589;
 wire m590;
 wire m591;
 wire m592;
 wire m593;
 wire m594;
 wire m595;
 wire m596;
 wire m597;
 wire m598;
 wire m599;
 wire m600;
 wire m601;
 wire m602;
 wire m603;
 wire m604;
 wire m605;
 wire m606;
 wire m607;
 wire m608;
 wire m609;
 wire m610;
 wire m611;
 wire m612;
 wire m613;
 wire m614;
 wire m615;
 wire m616;
 wire m617;
 wire m618;
 wire m619;
 wire m620;
 wire m621;
 wire m622;
 wire m623;
 wire m624;
 wire m625;
 wire m626;
 wire m627;
 wire m628;
 wire m629;
 wire m630;
 wire m631;
 wire m632;
 wire m633;
 wire m634;
 wire m635;
 wire m636;
 wire m637;
 wire m638;
 wire m639;
 wire m640;
 wire m641;
 wire m642;
 wire m643;
 wire m644;
 wire m645;
 wire m646;
 wire m647;
 wire m648;
 wire m649;
 wire m650;
 wire m651;
 wire m652;
 wire m653;
 wire m654;
 wire m655;
 wire m656;
 wire m657;
 wire m658;
 wire m659;
 wire m660;
 wire m661;
 wire m662;
 wire m663;
 wire m664;
 wire m665;
 wire m666;
 wire m667;
 wire m668;
 wire m669;
 wire m670;
 wire m671;
 wire m672;
 wire m673;
 wire m674;
 wire m675;
 wire m676;
 wire m677;
 wire m678;
 wire m679;
 wire m680;
 wire m681;
 wire m682;
 wire m683;
 wire m684;
 wire m685;
 wire m686;
 wire m687;
 wire m688;
 wire m689;
 wire m690;
 wire m691;
 wire m692;
 wire m693;
 wire m694;
 wire m695;
 wire m696;
 wire m697;
 wire m698;
 wire m699;
 wire m700;
 wire m701;
 wire m702;
 wire m703;
 wire m704;
 wire m705;
 wire m706;
 wire m707;
 wire m708;
 wire m709;
 wire m710;
 wire m711;
 wire m712;
 wire m713;
 wire m714;
 wire m715;
 wire m716;
 wire m717;
 wire m718;
 wire m719;
 wire m720;
 wire m721;
 wire m722;
 wire m723;
 wire m724;
 wire m725;
 wire m726;
 wire m727;
 wire m728;
 wire m729;
 wire m730;
 wire m731;
 wire m732;
 wire m733;
 wire m734;
 wire m735;
 wire m736;
 wire m737;
 wire m738;
 wire m739;
 wire m740;
 wire m741;
 wire m742;
 wire m743;
 wire m744;
 wire m745;
 wire m746;
 wire m747;
 wire m748;
 wire m749;
 wire m750;
 wire m751;
 wire m752;
 wire m753;
 wire m754;
 wire m755;
 wire m756;
 wire m757;
 wire m758;
 wire m759;
 wire m760;
 wire m761;
 wire m762;
 wire m763;
 wire m764;
 wire m765;
 wire m766;
 wire m767;
 wire m768;
 wire m769;
 wire m770;
 wire m771;
 wire m772;
 wire m773;
 wire m774;
 wire m775;
 wire m776;
 wire m777;
 wire m778;
 wire m779;
 wire m780;
 wire m781;
 wire m782;
 wire m783;
 wire m784;
 wire m785;
 wire m786;
 wire m787;
 wire m788;
 wire m789;
 wire m790;
 wire m791;
 wire m792;
 wire m793;
 wire m794;
 wire m795;
 wire m796;
 wire m797;
 wire m798;
 wire m799;
 wire m800;
 wire m801;
 wire m802;
 wire m803;
 wire m804;
 wire m805;
 wire m806;
 wire m807;
 wire m808;
 wire m809;
 wire m810;
 wire m811;
 wire m812;
 wire m813;
 wire m814;
 wire m815;
 wire m816;
 wire m817;
 wire m818;
 wire m819;
 wire m820;
 wire m821;
 wire m822;
 wire m823;
 wire m824;
 wire m825;
 wire m826;
 wire m827;
 wire m828;
 wire m829;
 wire m830;
 wire m831;
 wire m832;
 wire m833;
 wire m834;
 wire m835;
 wire m836;
 wire m837;
 wire m838;
 wire m839;
 wire m840;
 wire m841;
 wire m842;
 wire m843;
 wire m844;
 wire m845;
 wire m846;
 wire m847;
 wire m848;
 wire m849;
 wire m850;
 wire m851;
 wire m852;
 wire m853;
 wire m854;
 wire m855;
 wire m856;
 wire m857;
 wire m858;
 wire m859;
 wire m860;
 wire m861;
 wire m862;
 wire m863;
 wire m864;
 wire m865;
 wire m866;
 wire m867;
 wire m868;
 wire m869;
 wire m870;
 wire m871;
 wire m872;
 wire m873;
 wire m874;
 wire m875;
 wire m876;
 wire m877;
 wire m878;
 wire m879;
 wire m880;
 wire m881;
 wire m882;
 wire m883;
 wire m884;
 wire m885;
 wire m886;
 wire m887;
 wire m888;
 wire m889;
 wire m890;
 wire m891;
 wire m892;
 wire m893;
 wire m894;
 wire m895;
 wire m896;
 wire m897;
 wire m898;
 wire m899;
 wire m900;
 wire m901;
 wire m902;
 wire m903;
 wire m904;
 wire m905;
 wire m906;
 wire m907;
 wire m908;
 wire m909;
 wire m910;
 wire m911;
 wire m912;
 wire m913;
 wire m914;
 wire m915;
 wire m916;
 wire m917;
 wire m918;
 wire m919;
 wire m920;
 wire m921;
 wire m922;
 wire m923;
 wire m924;
 wire m925;
 wire m926;
 wire m927;
 wire m928;
 wire m929;
 wire m930;
 wire m931;
 wire m932;
 wire m933;
 wire m934;
 wire m935;
 wire m936;
 wire m937;
 wire m938;
 wire m939;
 wire m940;
 wire m941;
 wire m942;
 wire m943;
 wire m944;
 wire m945;
 wire m946;
 wire m947;
 wire m948;
 wire m949;
 wire m950;
 wire m951;
 wire m952;
 wire m953;
 wire m954;
 wire m955;
 wire m956;
 wire m957;
 wire m958;
 wire m959;
 wire m960;
 wire m961;
 wire m962;
 wire m963;
 wire m964;
 wire m965;
 wire m966;
 wire m967;
 wire m968;
 wire m969;
 wire m970;
 wire m971;
 wire m972;
 wire m973;
 wire m974;
 wire m975;
 wire m976;
 wire m977;
 wire m978;
 wire m979;
 wire m980;
 wire m981;
 wire m982;
 wire m983;
 wire m984;
 wire m985;
 wire m986;
 wire m987;
 wire m988;
 wire m989;
 wire m990;
 wire m991;
 wire m992;
 wire m993;
 wire m994;
 wire m995;
 wire m996;
 wire m997;
 wire m998;
 wire m999;
 wire m1000;
 wire m1001;
 wire m1002;
 wire m1003;
 wire m1004;
 wire m1005;
 wire m1006;
 wire m1007;
 wire m1008;
 wire m1009;
 wire m1010;
 wire m1011;
 wire m1012;
 wire m1013;
 wire m1014;
 wire m1015;
 wire m1016;
 wire m1017;
 wire m1018;
 wire m1019;
 wire m1020;
 wire m1021;
 wire m1022;
 wire m1023;
 wire m1024;
 wire m1025;
 wire m1026;
 wire m1027;
 wire m1028;
 wire m1029;
 wire m1030;
 wire m1031;
 wire m1032;
 wire m1033;
 wire m1034;
 wire m1035;
 wire m1036;
 wire m1037;
 wire m1038;
 wire m1039;
 wire m1040;
 wire m1041;
 wire m1042;
 wire m1043;
 wire m1044;
 wire m1045;
 wire m1046;
 wire m1047;
 wire m1048;
 wire m1049;
 wire m1050;
 wire m1051;
 wire m1052;
 wire m1053;
 wire m1054;
 wire m1055;
 wire m1056;
 wire m1057;
 wire m1058;
 wire m1059;
 wire m1060;
 wire m1061;
 wire m1062;
 wire m1063;
 wire m1064;
 wire m1065;
 wire m1066;
 wire m1067;
 wire m1068;
 wire m1069;
 wire m1070;
 wire m1071;
 wire m1072;
 wire m1073;
 wire m1074;
 wire m1075;
 wire m1076;
 wire m1077;
 wire m1078;
 wire m1079;
 wire m1080;
 wire m1081;
 wire m1082;
 wire m1083;
 wire m1084;
 wire m1085;
 wire m1086;
 wire m1087;
 wire m1088;
 wire m1089;
 wire m1090;
 wire m1091;
 wire m1092;
 wire m1093;
 wire m1094;
 wire m1095;
 wire m1096;
 wire m1097;
 wire m1098;
 wire m1099;
 wire m1100;
 wire m1101;
 wire m1102;
 wire m1103;
 wire m1104;
 wire m1105;
 wire m1106;
 wire m1107;
 wire m1108;
 wire m1109;
 wire m1110;
 wire m1111;
 wire m1112;
 wire m1113;
 wire m1114;
 wire m1115;
 wire m1116;
 wire m1117;
 wire m1118;
 wire m1119;
 wire m1120;
 wire m1121;
 wire m1122;
 wire m1123;
 wire m1124;
 wire m1125;
 wire m1126;
 wire m1127;
 wire m1128;
 wire m1129;
 wire m1130;
 wire m1131;
 wire m1132;
 wire m1133;
 wire m1134;
 wire m1135;
 wire m1136;
 wire m1137;
 wire m1138;
 wire m1139;
 wire m1140;
 wire m1141;
 wire m1142;
 wire m1143;
 wire m1144;
 wire m1145;
 wire m1146;
 wire m1147;
 wire m1148;
 wire m1149;
 wire m1150;
 wire m1151;
 wire m1152;
 wire m1153;
 wire m1154;
 wire m1155;
 wire m1156;
 wire m1157;
 wire m1158;
 wire m1159;
 wire m1160;
 wire m1161;
 wire m1162;
 wire m1163;
 wire m1164;
 wire m1165;
 wire m1166;
 wire m1167;
 wire m1168;
 wire m1169;
 wire m1170;
 wire m1171;
 wire m1172;
 wire m1173;
 wire m1174;
 wire m1175;
 wire m1176;
 wire m1177;
 wire m1178;
 wire m1179;
 wire m1180;
 wire m1181;
 wire m1182;
 wire m1183;
 wire m1184;
 wire m1185;
 wire m1186;
 wire m1187;
 wire m1188;
 wire m1189;
 wire m1190;
 wire m1191;
 wire m1192;
 wire m1193;
 wire m1194;
 wire m1195;
 wire m1196;
 wire m1197;
 wire m1198;
 wire m1199;
 wire m1200;
 wire m1201;
 m_12 inst_1(.i1(i12[1]),
            .i2(m6),
            .i3(m7),
            .o1(m158));
 m_12 inst_2(.i1(i12[0]),
            .i2(m6),
            .i3(m176),
            .o1(m1461));
 m_12 inst_3(.i1(m1),
            .i2(m1461),
            .i3(m5),
            .o1(o1[0]));
 m_8 inst_4(.i1(m2),
           .i2(m13),
           .o1(m1));
 m_14 inst_5(.i1(m3),
            .i2(m4),
            .i3(m228),
            .o1(m2));
 m_8 inst_6(.i1(i7[2]),
           .i2(i7[3]),
           .o1(m3));
 m_8 inst_7(.i1(i7[0]),
           .i2(i7[1]),
           .o1(m4));
 m_19 inst_8(.i1(i8[0]),
            .i2(m179),
            .i3(m166),
            .i4(i6[0]),
            .o1(m5));
 m_10 inst_9(.i1(i3[1]),
            .i2(i3[0]),
            .o1(m6));
 m_12 inst_10(.i1(m8),
             .i2(m9),
             .i3(m65),
             .o1(m7));
 m_12 inst_11(.i1(m10),
             .i2(m9),
             .i3(m11),
             .o1(m13));
 m_8 inst_12(.i1(m1322),
            .i2(m12),
            .o1(m11));
 m_14 inst_13(.i1(m64),
             .i2(m67),
             .i3(m14),
             .o1(m12));
 m_12 inst_14(.i1(m14),
             .i2(m15),
             .i3(m63),
             .o1(m9));
 m_5 inst_15(.i1(m16),
            .o1(m15));
 m_2 inst_16(.i1(i7[2]),
            .i2(i7[6]),
            .i3(m228),
            .o1(m16));
 m_10 inst_17(.i1(m14),
             .i2(m15),
             .o1(m17));
 m_12 inst_18(.i1(m14),
             .i2(m18),
             .i3(m17),
             .o1(m61));
 m_2 inst_19(.i1(m18),
            .i2(m19),
            .i3(m14),
            .o1(m59));
 m_2 inst_20(.i1(m19),
            .i2(m20),
            .i3(m14),
            .o1(m57));
 m_2 inst_21(.i1(m20),
            .i2(m21),
            .i3(m14),
            .o1(m55));
 m_2 inst_22(.i1(m21),
            .i2(m22),
            .i3(m14),
            .o1(m53));
 m_2 inst_23(.i1(m22),
            .i2(m23),
            .i3(m14),
            .o1(m51));
 m_2 inst_24(.i1(m23),
            .i2(m24),
            .i3(m14),
            .o1(m49));
 m_2 inst_25(.i1(m24),
            .i2(m25),
            .i3(m14),
            .o1(m47));
 m_2 inst_26(.i1(m25),
            .i2(m26),
            .i3(m14),
            .o1(m45));
 m_2 inst_27(.i1(m26),
            .i2(m27),
            .i3(m14),
            .o1(m42));
 m_2 inst_28(.i1(m27),
            .i2(m28),
            .i3(m14),
            .o1(m34));
 m_14 inst_29(.i1(m29),
             .i2(m28),
             .i3(m32),
             .o1(m82));
 m_8 inst_30(.i1(m30),
            .i2(m29),
            .o1(m10));
 m_5 inst_31(.i1(m33),
            .o1(m30));
 m_8 inst_32(.i1(m30),
            .i2(m31),
            .o1(m14));
 m_8 inst_33(.i1(m31),
            .i2(m79),
            .o1(m29));
 m_12 inst_34(.i1(m33),
             .i2(m31),
             .i3(m175),
             .o1(m32));
 m_14 inst_35(.i1(i7[27]),
             .i2(m228),
             .i3(i7[31]),
             .o1(m33));
 m_14 inst_36(.i1(i7[24]),
             .i2(m228),
             .i3(i7[28]),
             .o1(m28));
 m_8 inst_37(.i1(m8),
            .i2(m34),
            .o1(m35));
 m_8 inst_38(.i1(m10),
            .i2(m34),
            .o1(m92));
 m_12 inst_39(.i1(m35),
             .i2(m81),
             .i3(m36),
             .o1(m37));
 m_14 inst_40(.i1(i14),
             .i2(i6[23]),
             .i3(m179),
             .o1(m36));
 m_12 inst_41(.i1(i17),
             .i2(i8[23]),
             .i3(m37),
             .o1(m38));
 m_5 inst_42(.i1(m38),
            .o1(o1[23]));
 m_12 inst_43(.i1(i7[22]),
             .i2(m212),
             .i3(m39),
             .o1(m27));
 m_10 inst_44(.i1(m40),
             .i2(m212),
             .o1(m39));
 m_5 inst_45(.i1(i7[26]),
            .o1(m40));
 m_12 inst_46(.i1(m40),
             .i2(m212),
             .i3(m41),
             .o1(m31));
 m_5 inst_47(.i1(i7[30]),
            .o1(m41));
 m_8 inst_48(.i1(m10),
            .i2(m42),
            .o1(m43));
 m_12 inst_49(.i1(m8),
             .i2(m42),
             .i3(m175),
             .o1(m44));
 m_2 inst_50(.i1(i7[20]),
            .i2(i7[24]),
            .i3(m228),
            .o1(m26));
 m_12 inst_51(.i1(m8),
             .i2(m45),
             .i3(m175),
             .o1(m46));
 m_12 inst_52(.i1(m10),
             .i2(m45),
             .i3(m175),
             .o1(m107));
 m_2 inst_53(.i1(i7[18]),
            .i2(i7[22]),
            .i3(m228),
            .o1(m25));
 m_8 inst_54(.i1(m8),
            .i2(m47),
            .o1(m48));
 m_12 inst_55(.i1(m10),
             .i2(m47),
             .i3(m176),
             .o1(m115));
 m_2 inst_56(.i1(i7[16]),
            .i2(i7[20]),
            .i3(m228),
            .o1(m24));
 m_8 inst_57(.i1(m8),
            .i2(m49),
            .o1(m50));
 m_12 inst_58(.i1(m10),
             .i2(m49),
             .i3(m176),
             .o1(m121));
 m_2 inst_59(.i1(i7[14]),
            .i2(i7[18]),
            .i3(m228),
            .o1(m23));
 m_8 inst_60(.i1(m8),
            .i2(m51),
            .o1(m52));
 m_12 inst_61(.i1(m10),
             .i2(m51),
             .i3(m176),
             .o1(m127));
 m_2 inst_62(.i1(i7[12]),
            .i2(i7[16]),
            .i3(m228),
            .o1(m22));
 m_8 inst_63(.i1(m8),
            .i2(m53),
            .o1(m54));
 m_12 inst_64(.i1(m10),
             .i2(m53),
             .i3(m176),
             .o1(m133));
 m_2 inst_65(.i1(i7[10]),
            .i2(i7[14]),
            .i3(m228),
            .o1(m21));
 m_8 inst_66(.i1(m8),
            .i2(m55),
            .o1(m56));
 m_12 inst_67(.i1(m10),
             .i2(m55),
             .i3(m176),
             .o1(m139));
 m_2 inst_68(.i1(i7[8]),
            .i2(i7[12]),
            .i3(m228),
            .o1(m20));
 m_8 inst_69(.i1(m8),
            .i2(m57),
            .o1(m58));
 m_12 inst_70(.i1(m10),
             .i2(m57),
             .i3(m176),
             .o1(m145));
 m_2 inst_71(.i1(i7[6]),
            .i2(i7[10]),
            .i3(m228),
            .o1(m19));
 m_8 inst_72(.i1(m8),
            .i2(m59),
            .o1(m60));
 m_12 inst_73(.i1(m10),
             .i2(m59),
             .i3(m176),
             .o1(m151));
 m_2 inst_74(.i1(i7[4]),
            .i2(i7[8]),
            .i3(m228),
            .o1(m18));
 m_8 inst_75(.i1(m8),
            .i2(m61),
            .o1(m62));
 m_10 inst_76(.i1(m14),
             .i2(m64),
             .o1(m63));
 m_2 inst_77(.i1(i7[0]),
            .i2(i7[4]),
            .i3(m228),
            .o1(m64));
 m_14 inst_78(.i1(m8),
             .i2(m66),
             .i3(m1322),
             .o1(m65));
 m_2 inst_79(.i1(m67),
            .i2(m68),
            .i3(m14),
            .o1(m66));
 m_2 inst_80(.i1(i7[1]),
            .i2(i7[5]),
            .i3(m228),
            .o1(m67));
 m_2 inst_81(.i1(m68),
            .i2(m69),
            .i3(m14),
            .o1(m149));
 m_2 inst_82(.i1(m69),
            .i2(m70),
            .i3(m14),
            .o1(m143));
 m_2 inst_83(.i1(m70),
            .i2(m71),
            .i3(m14),
            .o1(m137));
 m_2 inst_84(.i1(m71),
            .i2(m72),
            .i3(m14),
            .o1(m131));
 m_2 inst_85(.i1(m72),
            .i2(m73),
            .i3(m14),
            .o1(m125));
 m_2 inst_86(.i1(m73),
            .i2(m74),
            .i3(m14),
            .o1(m119));
 m_2 inst_87(.i1(m74),
            .i2(m75),
            .i3(m14),
            .o1(m113));
 m_2 inst_88(.i1(m75),
            .i2(m76),
            .i3(m14),
            .o1(m105));
 m_2 inst_89(.i1(m76),
            .i2(m77),
            .i3(m14),
            .o1(m96));
 m_2 inst_90(.i1(m77),
            .i2(m78),
            .i3(m14),
            .o1(m86));
 m_2 inst_91(.i1(m78),
            .i2(m79),
            .i3(m14),
            .o1(m80));
 m_14 inst_92(.i1(i7[25]),
             .i2(m228),
             .i3(i7[29]),
             .o1(m79));
 m_12 inst_93(.i1(m31),
             .i2(m79),
             .i3(m33),
             .o1(m8));
 m_12 inst_94(.i1(m8),
             .i2(m80),
             .i3(m82),
             .o1(m83));
 m_12 inst_95(.i1(m10),
             .i2(m80),
             .i3(m175),
             .o1(m81));
 m_14 inst_96(.i1(m83),
             .i2(m84),
             .i3(m85),
             .o1(o1[24]));
 m_12 inst_97(.i1(m179),
             .i2(i6[24]),
             .i3(m159),
             .o1(m84));
 m_8 inst_98(.i1(i17),
            .i2(i8[24]),
            .o1(m85));
 m_2 inst_99(.i1(i7[27]),
            .i2(i7[23]),
            .i3(m212),
            .o1(m78));
 m_8 inst_100(.i1(m10),
             .i2(m86),
             .o1(m87));
 m_12 inst_101(.i1(m87),
              .i2(m44),
              .i3(m88),
              .o1(m89));
 m_14 inst_102(.i1(i14),
              .i2(i6[21]),
              .i3(m179),
              .o1(m88));
 m_12 inst_103(.i1(i17),
              .i2(i8[21]),
              .i3(m89),
              .o1(m90));
 m_5 inst_104(.i1(m90),
             .o1(o1[21]));
 m_12 inst_105(.i1(m8),
              .i2(m86),
              .i3(m175),
              .o1(m91));
 m_12 inst_106(.i1(m92),
              .i2(m91),
              .i3(m93),
              .o1(m94));
 m_14 inst_107(.i1(i14),
              .i2(i6[22]),
              .i3(m179),
              .o1(m93));
 m_12 inst_108(.i1(i17),
              .i2(i8[22]),
              .i3(m94),
              .o1(m95));
 m_5 inst_109(.i1(m95),
             .o1(o1[22]));
 m_2 inst_110(.i1(i7[25]),
             .i2(i7[21]),
             .i3(m212),
             .o1(m77));
 m_8 inst_111(.i1(m10),
             .i2(m96),
             .o1(m97));
 m_12 inst_112(.i1(m97),
              .i2(m46),
              .i3(m98),
              .o1(m99));
 m_14 inst_113(.i1(i14),
              .i2(i6[19]),
              .i3(m179),
              .o1(m98));
 m_12 inst_114(.i1(i17),
              .i2(i8[19]),
              .i3(m99),
              .o1(m100));
 m_5 inst_115(.i1(m100),
             .o1(o1[19]));
 m_12 inst_116(.i1(m8),
              .i2(m96),
              .i3(m175),
              .o1(m101));
 m_12 inst_117(.i1(m43),
              .i2(m101),
              .i3(m102),
              .o1(m103));
 m_14 inst_118(.i1(i14),
              .i2(i6[20]),
              .i3(m179),
              .o1(m102));
 m_12 inst_119(.i1(i17),
              .i2(i8[20]),
              .i3(m103),
              .o1(m104));
 m_5 inst_120(.i1(m104),
             .o1(o1[20]));
 m_2 inst_121(.i1(i7[19]),
             .i2(i7[23]),
             .i3(m228),
             .o1(m76));
 m_8 inst_122(.i1(m8),
             .i2(m105),
             .o1(m106));
 m_12 inst_123(.i1(m106),
              .i2(m107),
              .i3(m108),
              .o1(m109));
 m_14 inst_124(.i1(i14),
              .i2(i6[18]),
              .i3(m179),
              .o1(m108));
 m_12 inst_125(.i1(i17),
              .i2(i8[18]),
              .i3(m109),
              .o1(m110));
 m_5 inst_126(.i1(m110),
             .o1(o1[18]));
 m_12 inst_127(.i1(m10),
              .i2(m105),
              .i3(m176),
              .o1(m111));
 m_12 inst_128(.i1(m48),
              .i2(m111),
              .i3(m112),
              .o1(o1[17]));
 m_19 inst_129(.i1(m179),
              .i2(i8[17]),
              .i3(m166),
              .i4(i6[17]),
              .o1(m112));
 m_2 inst_130(.i1(i7[17]),
             .i2(i7[21]),
             .i3(m228),
             .o1(m75));
 m_8 inst_131(.i1(m8),
             .i2(m113),
             .o1(m114));
 m_12 inst_132(.i1(m114),
              .i2(m115),
              .i3(m116),
              .o1(o1[16]));
 m_19 inst_133(.i1(m179),
              .i2(i8[16]),
              .i3(m166),
              .i4(i6[16]),
              .o1(m116));
 m_12 inst_134(.i1(m10),
              .i2(m113),
              .i3(m176),
              .o1(m117));
 m_12 inst_135(.i1(m50),
              .i2(m117),
              .i3(m118),
              .o1(o1[15]));
 m_19 inst_136(.i1(m179),
              .i2(i8[15]),
              .i3(m166),
              .i4(i6[15]),
              .o1(m118));
 m_2 inst_137(.i1(i7[15]),
             .i2(i7[19]),
             .i3(m228),
             .o1(m74));
 m_8 inst_138(.i1(m8),
             .i2(m119),
             .o1(m120));
 m_12 inst_139(.i1(m120),
              .i2(m121),
              .i3(m122),
              .o1(o1[14]));
 m_19 inst_140(.i1(m179),
              .i2(i8[14]),
              .i3(m166),
              .i4(i6[14]),
              .o1(m122));
 m_12 inst_141(.i1(m10),
              .i2(m119),
              .i3(m176),
              .o1(m123));
 m_12 inst_142(.i1(m52),
              .i2(m123),
              .i3(m124),
              .o1(o1[13]));
 m_19 inst_143(.i1(m179),
              .i2(i8[13]),
              .i3(m166),
              .i4(i6[13]),
              .o1(m124));
 m_2 inst_144(.i1(i7[13]),
             .i2(i7[17]),
             .i3(m228),
             .o1(m73));
 m_8 inst_145(.i1(m8),
             .i2(m125),
             .o1(m126));
 m_12 inst_146(.i1(m126),
              .i2(m127),
              .i3(m128),
              .o1(o1[12]));
 m_19 inst_147(.i1(m179),
              .i2(i8[12]),
              .i3(m166),
              .i4(i6[12]),
              .o1(m128));
 m_12 inst_148(.i1(m10),
              .i2(m125),
              .i3(m176),
              .o1(m129));
 m_12 inst_149(.i1(m54),
              .i2(m129),
              .i3(m130),
              .o1(o1[11]));
 m_19 inst_150(.i1(m179),
              .i2(i8[11]),
              .i3(m166),
              .i4(i6[11]),
              .o1(m130));
 m_2 inst_151(.i1(i7[11]),
             .i2(i7[15]),
             .i3(m228),
             .o1(m72));
 m_8 inst_152(.i1(m8),
             .i2(m131),
             .o1(m132));
 m_12 inst_153(.i1(m132),
              .i2(m133),
              .i3(m134),
              .o1(o1[10]));
 m_19 inst_154(.i1(m179),
              .i2(i8[10]),
              .i3(m166),
              .i4(i6[10]),
              .o1(m134));
 m_12 inst_155(.i1(m10),
              .i2(m131),
              .i3(m176),
              .o1(m135));
 m_12 inst_156(.i1(m56),
              .i2(m135),
              .i3(m136),
              .o1(o1[9]));
 m_19 inst_157(.i1(m179),
              .i2(i8[9]),
              .i3(m166),
              .i4(i6[9]),
              .o1(m136));
 m_2 inst_158(.i1(i7[9]),
             .i2(i7[13]),
             .i3(m228),
             .o1(m71));
 m_8 inst_159(.i1(m8),
             .i2(m137),
             .o1(m138));
 m_12 inst_160(.i1(m138),
              .i2(m139),
              .i3(m140),
              .o1(o1[8]));
 m_19 inst_161(.i1(m179),
              .i2(i8[8]),
              .i3(m166),
              .i4(i6[8]),
              .o1(m140));
 m_12 inst_162(.i1(m10),
              .i2(m137),
              .i3(m176),
              .o1(m141));
 m_12 inst_163(.i1(m58),
              .i2(m141),
              .i3(m142),
              .o1(o1[7]));
 m_19 inst_164(.i1(m179),
              .i2(i8[7]),
              .i3(m166),
              .i4(i6[7]),
              .o1(m142));
 m_2 inst_165(.i1(i7[7]),
             .i2(i7[11]),
             .i3(m228),
             .o1(m70));
 m_8 inst_166(.i1(m8),
             .i2(m143),
             .o1(m144));
 m_12 inst_167(.i1(m144),
              .i2(m145),
              .i3(m146),
              .o1(o1[6]));
 m_19 inst_168(.i1(m179),
              .i2(i8[6]),
              .i3(m166),
              .i4(i6[6]),
              .o1(m146));
 m_12 inst_169(.i1(m10),
              .i2(m143),
              .i3(m176),
              .o1(m147));
 m_12 inst_170(.i1(m60),
              .i2(m147),
              .i3(m148),
              .o1(o1[5]));
 m_19 inst_171(.i1(m179),
              .i2(i8[5]),
              .i3(m166),
              .i4(i6[5]),
              .o1(m148));
 m_2 inst_172(.i1(i7[5]),
             .i2(i7[9]),
             .i3(m228),
             .o1(m69));
 m_8 inst_173(.i1(m8),
             .i2(m149),
             .o1(m150));
 m_12 inst_174(.i1(m150),
              .i2(m151),
              .i3(m152),
              .o1(o1[4]));
 m_19 inst_175(.i1(m179),
              .i2(i8[4]),
              .i3(m166),
              .i4(i6[4]),
              .o1(m152));
 m_12 inst_176(.i1(m10),
              .i2(m149),
              .i3(m176),
              .o1(m153));
 m_12 inst_177(.i1(m62),
              .i2(m153),
              .i3(m154),
              .o1(o1[3]));
 m_19 inst_178(.i1(m179),
              .i2(i8[3]),
              .i3(m166),
              .i4(i6[3]),
              .o1(m154));
 m_2 inst_179(.i1(i7[3]),
             .i2(i7[7]),
             .i3(m228),
             .o1(m68));
 m_8 inst_180(.i1(m8),
             .i2(m66),
             .o1(m155));
 m_12 inst_181(.i1(m155),
              .i2(m156),
              .i3(m157),
              .o1(o1[2]));
 m_12 inst_182(.i1(m10),
              .i2(m61),
              .i3(m176),
              .o1(m156));
 m_19 inst_183(.i1(m179),
              .i2(i8[2]),
              .i3(m166),
              .i4(i6[2]),
              .o1(m157));
 m_12 inst_184(.i1(m159),
              .i2(m158),
              .i3(m165),
              .o1(o1[1]));
 m_14 inst_185(.i1(i15[9]),
              .i2(m169),
              .i3(m159),
              .o1(m160));
 m_12 inst_186(.i1(i15[9]),
              .i2(m169),
              .i3(m160),
              .o1(m161));
 m_12 inst_187(.i1(i17),
              .i2(m162),
              .i3(m161),
              .o1(o1[34]));
 m_5 inst_188(.i1(i8[34]),
             .o1(m162));
 m_10 inst_189(.i1(m175),
              .i2(i17),
              .o1(m159));
 m_12 inst_190(.i1(m159),
              .i2(m163),
              .i3(m164),
              .o1(o1[25]));
 m_20 inst_191(.i1(i15[0]),
              .i2(m8),
              .o1(m163));
 m_19 inst_192(.i1(m179),
              .i2(i8[25]),
              .i3(m166),
              .i4(i6[25]),
              .o1(m164));
 m_19 inst_193(.i1(m179),
              .i2(i8[1]),
              .i3(m166),
              .i4(i6[1]),
              .o1(m165));
 m_8 inst_194(.i1(i14),
             .i2(i13),
             .o1(m167));
 m_12 inst_195(.i1(i15[8]),
              .i2(m168),
              .i3(m167),
              .o1(m170));
 m_8 inst_196(.i1(i15[8]),
             .i2(m168),
             .o1(m169));
 m_12 inst_197(.i1(m171),
              .i2(m170),
              .i3(i17),
              .o1(m172));
 m_15 inst_198(.i1(i15[8]),
              .i2(m168),
              .o1(m171));
 m_12 inst_199(.i1(m173),
              .i2(m172),
              .i3(m174),
              .o1(o1[33]));
 m_8 inst_200(.i1(m175),
             .i2(i6[33]),
             .o1(m173));
 m_10 inst_201(.i1(m179),
              .i2(i8[33]),
              .o1(m174));
 m_5 inst_202(.i1(i14),
             .o1(m175));
 m_8 inst_203(.i1(m175),
             .i2(m179),
             .o1(m166));
 m_8 inst_204(.i1(i14),
             .i2(m179),
             .o1(m176));
 m_10 inst_205(.i1(i17),
              .i2(i16),
              .o1(m177));
 m_12 inst_206(.i1(i17),
              .i2(m178),
              .i3(m177),
              .o1(o1[35]));
 m_5 inst_207(.i1(i8[35]),
             .o1(m178));
 m_5 inst_208(.i1(i17),
             .o1(m179));
 m_10 inst_209(.i1(i17),
              .i2(i19),
              .o1(m180));
 m_12 inst_210(.i1(i17),
              .i2(m181),
              .i3(m180),
              .o1(o1[36]));
 m_5 inst_211(.i1(i8[36]),
             .o1(m181));
 m_12 inst_212(.i1(m182),
              .i2(m183),
              .i3(i2[0]),
              .o1(m184));
 m_8 inst_213(.i1(m182),
             .i2(m183),
             .o1(m1200));
 m_16 inst_214(.i1(m182),
              .i2(m183),
              .o1(m185));
 m_12 inst_215(.i1(m267),
              .i2(m185),
              .i3(m184),
              .o1(o20[23]));
 m_8 inst_216(.i1(i9[0]),
             .i2(m186),
             .o1(m187));
 m_5 inst_217(.i1(i15[3]),
             .o1(m186));
 m_8 inst_218(.i1(m187),
             .i2(m188),
             .o1(m189));
 m_12 inst_219(.i1(i9[1]),
              .i2(m190),
              .i3(m191),
              .o1(m192));
 m_5 inst_220(.i1(i15[4]),
             .o1(m190));
 m_12 inst_221(.i1(m187),
              .i2(m188),
              .i3(m207),
              .o1(m191));
 m_14 inst_222(.i1(i15[5]),
              .i2(m192),
              .i3(i14),
              .o1(m193));
 m_15 inst_223(.i1(m197),
              .i2(m193),
              .o1(m194));
 m_12 inst_224(.i1(m195),
              .i2(m194),
              .i3(m196),
              .o1(o1[30]));
 m_12 inst_225(.i1(m175),
              .i2(i6[30]),
              .i3(i17),
              .o1(m195));
 m_10 inst_226(.i1(m179),
              .i2(i8[30]),
              .o1(m196));
 m_16 inst_227(.i1(i15[5]),
              .i2(m192),
              .o1(m197));
 m_14 inst_228(.i1(i15[6]),
              .i2(m197),
              .i3(i14),
              .o1(m198));
 m_15 inst_229(.i1(m202),
              .i2(m198),
              .o1(m199));
 m_12 inst_230(.i1(m200),
              .i2(m199),
              .i3(m201),
              .o1(o1[31]));
 m_12 inst_231(.i1(m175),
              .i2(i6[31]),
              .i3(i17),
              .o1(m200));
 m_10 inst_232(.i1(m179),
              .i2(i8[31]),
              .o1(m201));
 m_16 inst_233(.i1(i15[6]),
              .i2(m197),
              .o1(m202));
 m_14 inst_234(.i1(i15[7]),
              .i2(m202),
              .i3(i14),
              .o1(m203));
 m_15 inst_235(.i1(m168),
              .i2(m203),
              .o1(m204));
 m_12 inst_236(.i1(m205),
              .i2(m204),
              .i3(m206),
              .o1(o1[32]));
 m_12 inst_237(.i1(m175),
              .i2(i6[32]),
              .i3(i17),
              .o1(m205));
 m_10 inst_238(.i1(m179),
              .i2(i8[32]),
              .o1(m206));
 m_16 inst_239(.i1(i15[7]),
              .i2(m202),
              .o1(m168));
 m_6 inst_240(.i1(i9[1]),
             .i2(i15[4]),
             .o1(m207));
 m_20 inst_241(.i1(m189),
              .i2(m207),
              .o1(m208));
 m_12 inst_242(.i1(m159),
              .i2(m208),
              .i3(m209),
              .o1(o1[29]));
 m_19 inst_243(.i1(m179),
              .i2(i8[29]),
              .i3(m166),
              .i4(i6[29]),
              .o1(m209));
 m_20 inst_244(.i1(i9[0]),
              .i2(i15[3]),
              .o1(m210));
 m_14 inst_245(.i1(m211),
              .i2(m215),
              .i3(m210),
              .o1(m188));
 m_10 inst_246(.i1(i15[2]),
              .i2(m212),
              .o1(m211));
 m_10 inst_247(.i1(m213),
              .i2(m214),
              .o1(m212));
 m_15 inst_248(.i1(m213),
              .i2(m214),
              .o1(m228));
 m_8 inst_249(.i1(i7[29]),
             .i2(i7[28]),
             .o1(m213));
 m_8 inst_250(.i1(i7[31]),
             .i2(i7[30]),
             .o1(m214));
 m_10 inst_251(.i1(m176),
              .i2(m215),
              .o1(m216));
 m_12 inst_252(.i1(m219),
              .i2(m216),
              .i3(m217),
              .o1(o1[27]));
 m_19 inst_253(.i1(m179),
              .i2(i8[27]),
              .i3(m166),
              .i4(i6[27]),
              .o1(m217));
 m_10 inst_254(.i1(m218),
              .i2(m227),
              .o1(m215));
 m_8 inst_255(.i1(m218),
             .i2(m227),
             .o1(m219));
 m_12 inst_256(.i1(m220),
              .i2(m14),
              .i3(m221),
              .o1(m218));
 m_5 inst_257(.i1(i15[1]),
             .o1(m220));
 m_12 inst_258(.i1(i15[0]),
              .i2(m8),
              .i3(m222),
              .o1(m221));
 m_15 inst_259(.i1(m223),
              .i2(m222),
              .o1(m224));
 m_16 inst_260(.i1(i15[0]),
              .i2(m8),
              .o1(m223));
 m_12 inst_261(.i1(m224),
              .i2(m226),
              .i3(m225),
              .o1(o1[26]));
 m_19 inst_262(.i1(m179),
              .i2(i8[26]),
              .i3(m166),
              .i4(i6[26]),
              .o1(m225));
 m_12 inst_263(.i1(m223),
              .i2(m222),
              .i3(m176),
              .o1(m226));
 m_6 inst_264(.i1(i15[1]),
             .i2(m14),
             .o1(m222));
 m_6 inst_265(.i1(i15[2]),
             .i2(m228),
             .o1(m227));
 m_13 inst_266(.i1(m211),
              .i2(m215),
              .i3(m210),
              .o1(m229));
 m_10 inst_267(.i1(m176),
              .i2(m229),
              .o1(m230));
 m_12 inst_268(.i1(m188),
              .i2(m230),
              .i3(m231),
              .o1(o1[28]));
 m_19 inst_269(.i1(m179),
              .i2(i8[28]),
              .i3(m166),
              .i4(i6[28]),
              .o1(m231));
 m_12 inst_270(.i1(m1454),
              .i2(m232),
              .i3(m233),
              .o1(o10));
 m_10 inst_271(.i1(m1454),
              .i2(o6[33]),
              .o1(m233));
 m_13 inst_272(.i1(m1454),
              .i2(m234),
              .i3(m299),
              .o1(o11));
 m_13 inst_273(.i1(m235),
              .i2(m238),
              .i3(m259),
              .o1(m234));
 m_8 inst_274(.i1(m236),
             .i2(m237),
             .o1(m235));
 m_5 inst_275(.i1(m239),
             .o1(m238));
 m_13 inst_276(.i1(m308),
              .i2(m238),
              .i3(m240),
              .o1(m241));
 m_10 inst_277(.i1(m241),
              .i2(m242),
              .o1(m243));
 m_13 inst_278(.i1(m241),
              .i2(m242),
              .i3(m252),
              .o1(m253));
 m_13 inst_279(.i1(m241),
              .i2(m242),
              .i3(m244),
              .o1(m248));
 m_19 inst_280(.i1(m245),
              .i2(m1198),
              .i3(m276),
              .i4(m247),
              .o1(m244));
 m_5 inst_281(.i1(i4[12]),
             .o1(m245));
 m_12 inst_282(.i1(m245),
              .i2(m185),
              .i3(m246),
              .o1(o20[13]));
 m_12 inst_283(.i1(m182),
              .i2(m183),
              .i3(i4[13]),
              .o1(m246));
 m_19 inst_284(.i1(m1454),
              .i2(i5[12]),
              .i3(m929),
              .i4(i4[12]),
              .o1(m247));
 m_12 inst_285(.i1(m257),
              .i2(m249),
              .i3(m248),
              .o1(m1012));
 m_17 inst_286(.i1(i4[11]),
              .i2(m314),
              .i3(m240),
              .i4(m250),
              .o1(m249));
 m_8 inst_287(.i1(m240),
             .i2(m250),
             .o1(m1156));
 m_12 inst_288(.i1(i3[1]),
              .i2(m786),
              .i3(m251),
              .o1(m250));
 m_10 inst_289(.i1(i4[11]),
              .i2(m929),
              .o1(m251));
 m_13 inst_290(.i1(m253),
              .i2(m258),
              .i3(m254),
              .o1(m965));
 m_12 inst_291(.i1(m255),
              .i2(m256),
              .i3(m244),
              .o1(m254));
 m_8 inst_292(.i1(m255),
             .i2(m256),
             .o1(m257));
 m_12 inst_293(.i1(m257),
              .i2(m258),
              .i3(m253),
              .o1(m999));
 m_17 inst_294(.i1(i4[13]),
              .i2(m314),
              .i3(m240),
              .i4(m1128),
              .o1(m258));
 m_13 inst_295(.i1(m259),
              .i2(m260),
              .i3(m266),
              .o1(m272));
 m_8 inst_296(.i1(m237),
             .i2(m261),
             .o1(m260));
 m_12 inst_297(.i1(i4[22]),
              .i2(m262),
              .i3(m1200),
              .o1(m261));
 m_5 inst_298(.i1(i5[22]),
             .o1(m262));
 m_12 inst_299(.i1(m262),
              .i2(m1200),
              .i3(m263),
              .o1(o21[22]));
 m_10 inst_300(.i1(i5[21]),
              .i2(m1200),
              .o1(m263));
 m_12 inst_301(.i1(m1195),
              .i2(m1196),
              .i3(m262),
              .o1(m264));
 m_12 inst_302(.i1(i4[22]),
              .i2(m1198),
              .i3(m264),
              .o1(m265));
 m_5 inst_303(.i1(m265),
             .o1(o17[22]));
 m_12 inst_304(.i1(m267),
              .i2(i5[22]),
              .i3(m268),
              .o1(m266));
 m_5 inst_305(.i1(i4[22]),
             .o1(m267));
 m_12 inst_306(.i1(m269),
              .i2(m270),
              .i3(m271),
              .o1(m268));
 m_12 inst_307(.i1(m853),
              .i2(i5[21]),
              .i3(m840),
              .o1(m271));
 m_5 inst_308(.i1(m272),
             .o1(m273));
 m_14 inst_309(.i1(m274),
              .i2(m273),
              .i3(m314),
              .o1(m1203));
 m_8 inst_310(.i1(m275),
             .i2(m239),
             .o1(m274));
 m_18 inst_311(.i1(m275),
              .i2(m239),
              .i3(m276),
              .o1(m255));
 m_12 inst_312(.i1(m1195),
              .i2(m1196),
              .i3(m1454),
              .o1(m276));
 m_12 inst_313(.i1(m314),
              .i2(m275),
              .i3(m295),
              .o1(m277));
 m_19 inst_314(.i1(i4[23]),
              .i2(i3[1]),
              .i3(m277),
              .i4(m278),
              .o1(m1293));
 m_8 inst_315(.i1(i3[1]),
             .i2(m185),
             .o1(m278));
 m_8 inst_316(.i1(m279),
             .i2(m289),
             .o1(m259));
 m_10 inst_317(.i1(m279),
              .i2(m289),
              .o1(m324));
 m_12 inst_318(.i1(m236),
              .i2(m279),
              .i3(m280),
              .o1(m287));
 m_14 inst_319(.i1(m281),
              .i2(m286),
              .i3(i3[1]),
              .o1(m280));
 m_19 inst_320(.i1(m1208),
              .i2(m282),
              .i3(m285),
              .i4(m281),
              .o1(m242));
 m_5 inst_321(.i1(m283),
             .o1(m282));
 m_12 inst_322(.i1(i4[27]),
              .i2(m1210),
              .i3(i3[1]),
              .o1(m283));
 m_10 inst_323(.i1(m1208),
              .i2(m282),
              .o1(m284));
 m_8 inst_324(.i1(i3[1]),
             .i2(m737),
             .o1(m285));
 m_6 inst_325(.i1(m706),
             .i2(m183),
             .o1(m286));
 m_12 inst_326(.i1(m703),
              .i2(m1454),
              .i3(m287),
              .o1(m938));
 m_6 inst_327(.i1(m288),
             .i2(m182),
             .o1(m279));
 m_6 inst_328(.i1(i4[24]),
             .i2(i5[24]),
             .o1(m288));
 m_15 inst_329(.i1(m692),
              .i2(m290),
              .o1(m289));
 m_13 inst_330(.i1(m291),
              .i2(m292),
              .i3(m294),
              .o1(m290));
 m_20 inst_331(.i1(i4[25]),
              .i2(i5[25]),
              .o1(m291));
 m_14 inst_332(.i1(m292),
              .i2(m294),
              .i3(m291),
              .o1(m293));
 m_10 inst_333(.i1(m703),
              .i2(i5[24]),
              .o1(m292));
 m_12 inst_334(.i1(m705),
              .i2(i5[23]),
              .i3(m288),
              .o1(m294));
 m_17 inst_335(.i1(m295),
              .i2(m712),
              .i3(m289),
              .i4(m236),
              .o1(m296));
 m_12 inst_336(.i1(i3[1]),
              .i2(m296),
              .i3(m297),
              .o1(m945));
 m_12 inst_337(.i1(m1215),
              .i2(m298),
              .i3(i3[1]),
              .o1(m297));
 m_8 inst_338(.i1(i4[25]),
             .i2(i4[24]),
             .o1(m298));
 m_12 inst_339(.i1(m300),
              .i2(m309),
              .i3(m313),
              .o1(m299));
 m_14 inst_340(.i1(m301),
              .i2(m302),
              .i3(m303),
              .o1(m300));
 m_10 inst_341(.i1(o17[30]),
              .i2(m312),
              .o1(m303));
 m_18 inst_342(.i1(m300),
              .i2(m309),
              .i3(m304),
              .o1(m308));
 m_12 inst_343(.i1(m310),
              .i2(m316),
              .i3(m305),
              .o1(m304));
 m_6 inst_344(.i1(m306),
             .i2(m746),
             .o1(m305));
 m_12 inst_345(.i1(i4[27]),
              .i2(m307),
              .i3(m661),
              .o1(m306));
 m_5 inst_346(.i1(i5[27]),
             .o1(m307));
 m_10 inst_347(.i1(i4[27]),
              .i2(m307),
              .o1(m657));
 m_12 inst_348(.i1(m1195),
              .i2(m1196),
              .i3(m308),
              .o1(m236));
 m_18 inst_349(.i1(m630),
              .i2(m310),
              .i3(m311),
              .o1(m309));
 m_15 inst_350(.i1(o17[30]),
              .i2(m312),
              .o1(m311));
 m_10 inst_351(.i1(i4[30]),
              .i2(i5[30]),
              .o1(m312));
 m_15 inst_352(.i1(m314),
              .i2(m315),
              .o1(m313));
 m_8 inst_353(.i1(m1195),
             .i2(m1196),
             .o1(m314));
 m_18 inst_354(.i1(m310),
              .i2(m316),
              .i3(m317),
              .o1(m315));
 m_13 inst_355(.i1(m318),
              .i2(m239),
              .i3(m323),
              .o1(m317));
 m_14 inst_356(.i1(m302),
              .i2(m319),
              .i3(m318),
              .o1(m320));
 m_13 inst_357(.i1(m645),
              .i2(m646),
              .i3(m647),
              .o1(m319));
 m_13 inst_358(.i1(m321),
              .i2(m322),
              .i3(m320),
              .o1(m275));
 m_12 inst_359(.i1(m630),
              .i2(m310),
              .i3(m311),
              .o1(m321));
 m_13 inst_360(.i1(m301),
              .i2(m302),
              .i3(m303),
              .o1(m322));
 m_20 inst_361(.i1(m306),
              .i2(m746),
              .o1(m318));
 m_8 inst_362(.i1(m324),
             .i2(m325),
             .o1(m323));
 m_12 inst_363(.i1(m182),
              .i2(m183),
              .i3(m237),
              .o1(m325));
 m_12 inst_364(.i1(i3[1]),
              .i2(m326),
              .i3(m330),
              .o1(o12));
 m_10 inst_365(.i1(m327),
              .i2(m328),
              .o1(m326));
 m_5 inst_366(.i1(i2[0]),
             .o1(m327));
 m_8 inst_367(.i1(m327),
             .i2(m185),
             .o1(o20[24]));
 m_5 inst_368(.i1(i2[1]),
             .o1(m328));
 m_8 inst_369(.i1(m328),
             .i2(m185),
             .o1(o21[24]));
 m_12 inst_370(.i1(m328),
              .i2(m1200),
              .i3(m329),
              .o1(o21[23]));
 m_10 inst_371(.i1(i5[22]),
              .i2(m1200),
              .o1(m329));
 m_13 inst_372(.i1(o19),
              .i2(m331),
              .i3(m526),
              .o1(m330));
 m_8 inst_373(.i1(m332),
             .i2(m395),
             .o1(m331));
 m_13 inst_374(.i1(m333),
              .i2(m358),
              .i3(m380),
              .o1(m332));
 m_12 inst_375(.i1(m620),
              .i2(m333),
              .i3(m334),
              .o1(m339));
 m_12 inst_376(.i1(m1454),
              .i2(m335),
              .i3(m572),
              .o1(m334));
 m_10 inst_377(.i1(m1454),
              .i2(m335),
              .o1(m624));
 m_20 inst_378(.i1(m336),
              .i2(m337),
              .o1(m335));
 m_12 inst_379(.i1(i4[31]),
              .i2(m698),
              .i3(m338),
              .o1(m337));
 m_14 inst_380(.i1(i4[26]),
              .i2(i4[31]),
              .i3(m1302),
              .o1(m338));
 m_5 inst_381(.i1(m339),
             .o1(m340));
 m_12 inst_382(.i1(m1454),
              .i2(m341),
              .i3(m607),
              .o1(m333));
 m_10 inst_383(.i1(m1454),
              .i2(m341),
              .o1(m342));
 m_12 inst_384(.i1(m1454),
              .i2(m343),
              .i3(m342),
              .o1(m627));
 m_12 inst_385(.i1(i3[1]),
              .i2(m343),
              .i3(m344),
              .o1(m357));
 m_10 inst_386(.i1(i3[1]),
              .i2(m345),
              .o1(m344));
 m_6 inst_387(.i1(i4[2]),
             .i2(m346),
             .o1(m345));
 m_12 inst_388(.i1(i4[0]),
              .i2(i4[1]),
              .i3(m1309),
              .o1(m346));
 m_6 inst_389(.i1(i4[6]),
             .i2(m347),
             .o1(m343));
 m_14 inst_390(.i1(m821),
              .i2(m393),
              .i3(m232),
              .o1(m347));
 m_20 inst_391(.i1(m348),
              .i2(m351),
              .o1(m341));
 m_10 inst_392(.i1(m348),
              .i2(m351),
              .o1(m349));
 m_13 inst_393(.i1(m348),
              .i2(m351),
              .i3(m350),
              .o1(m513));
 m_5 inst_394(.i1(m362),
             .o1(m350));
 m_6 inst_395(.i1(m614),
             .i2(m352),
             .o1(m351));
 m_12 inst_396(.i1(i1[1]),
              .i2(i1[0]),
              .i3(m791),
              .o1(m352));
 m_16 inst_397(.i1(o19),
              .i2(m333),
              .o1(m353));
 m_2 inst_398(.i1(m353),
             .i2(m354),
             .i3(o18),
             .o1(o5[18]));
 m_14 inst_399(.i1(o19),
              .i2(m357),
              .i3(m355),
              .o1(m354));
 m_12 inst_400(.i1(m605),
              .i2(m354),
              .i3(m340),
              .o1(o5[26]));
 m_2 inst_401(.i1(m356),
             .i2(m353),
             .i3(o18),
             .o1(o5[10]));
 m_10 inst_402(.i1(m620),
              .i2(m357),
              .o1(m356));
 m_8 inst_403(.i1(o18),
             .i2(m356),
             .o1(o5[2]));
 m_8 inst_404(.i1(m359),
             .i2(m377),
             .o1(m358));
 m_2 inst_405(.i1(m360),
             .i2(m364),
             .i3(m1454),
             .o1(m359));
 m_10 inst_406(.i1(m513),
              .i2(m361),
              .o1(m360));
 m_10 inst_407(.i1(m349),
              .i2(m362),
              .o1(m361));
 m_6 inst_408(.i1(m614),
             .i2(m363),
             .o1(m362));
 m_8 inst_409(.i1(i4[11]),
             .i2(m1261),
             .o1(m363));
 m_12 inst_410(.i1(i3[1]),
              .i2(m364),
              .i3(m365),
              .o1(m379));
 m_10 inst_411(.i1(i3[1]),
              .i2(m366),
              .o1(m365));
 m_6 inst_412(.i1(m367),
             .i2(m369),
             .o1(m366));
 m_5 inst_413(.i1(i4[3]),
             .o1(m367));
 m_12 inst_414(.i1(m367),
              .i2(m185),
              .i3(m368),
              .o1(o20[4]));
 m_12 inst_415(.i1(m182),
              .i2(m183),
              .i3(i4[4]),
              .o1(m368));
 m_14 inst_416(.i1(m879),
              .i2(m370),
              .i3(m232),
              .o1(m369));
 m_13 inst_417(.i1(m879),
              .i2(m367),
              .i3(m370),
              .o1(m392));
 m_8 inst_418(.i1(i4[1]),
             .i2(i4[2]),
             .o1(m370));
 m_20 inst_419(.i1(m371),
              .i2(m375),
              .o1(m364));
 m_10 inst_420(.i1(m1309),
              .i2(m372),
              .o1(m371));
 m_13 inst_421(.i1(m1309),
              .i2(m372),
              .i3(m452),
              .o1(m384));
 m_18 inst_422(.i1(i4[4]),
              .i2(m392),
              .i3(m373),
              .o1(m372));
 m_8 inst_423(.i1(i4[7]),
             .i2(m373),
             .o1(m374));
 m_10 inst_424(.i1(m393),
              .i2(m374),
              .o1(m1319));
 m_16 inst_425(.i1(i4[5]),
              .i2(i4[6]),
              .o1(m373));
 m_12 inst_426(.i1(m815),
              .i2(m1305),
              .i3(m376),
              .o1(m375));
 m_10 inst_427(.i1(m815),
              .i2(m1309),
              .o1(m376));
 m_16 inst_428(.i1(m378),
              .i2(m379),
              .o1(m377));
 m_10 inst_429(.i1(m620),
              .i2(m378),
              .o1(m483));
 m_10 inst_430(.i1(m620),
              .i2(m379),
              .o1(m500));
 m_8 inst_431(.i1(m381),
             .i2(m387),
             .o1(m380));
 m_10 inst_432(.i1(m620),
              .i2(m381),
              .o1(m482));
 m_12 inst_433(.i1(i3[1]),
              .i2(m512),
              .i3(m382),
              .o1(m381));
 m_10 inst_434(.i1(i3[1]),
              .i2(m383),
              .o1(m382));
 m_20 inst_435(.i1(m384),
              .i2(m385),
              .o1(m383));
 m_6 inst_436(.i1(m614),
             .i2(m386),
             .o1(m385));
 m_8 inst_437(.i1(i4[8]),
             .i2(m1261),
             .o1(m386));
 m_10 inst_438(.i1(m620),
              .i2(m387),
              .o1(m388));
 m_8 inst_439(.i1(o18),
             .i2(m388),
             .o1(o5[4]));
 m_12 inst_440(.i1(m1454),
              .i2(m389),
              .i3(m394),
              .o1(m387));
 m_12 inst_441(.i1(i3[1]),
              .i2(m389),
              .i3(m390),
              .o1(m378));
 m_10 inst_442(.i1(i4[0]),
              .i2(i3[1]),
              .o1(m390));
 m_6 inst_443(.i1(m887),
             .i2(m391),
             .o1(m389));
 m_10 inst_444(.i1(m392),
              .i2(m1309),
              .o1(m391));
 m_8 inst_445(.i1(i4[4]),
             .i2(m392),
             .o1(m393));
 m_10 inst_446(.i1(m1454),
              .i2(m383),
              .o1(m394));
 m_13 inst_447(.i1(m396),
              .i2(m509),
              .i3(m517),
              .o1(m395));
 m_8 inst_448(.i1(m397),
             .i2(m428),
             .o1(m396));
 m_8 inst_449(.i1(i3[1]),
             .i2(m398),
             .o1(m397));
 m_10 inst_450(.i1(i3[1]),
              .i2(m398),
              .o1(m399));
 m_14 inst_451(.i1(m399),
              .i2(m400),
              .i3(m407),
              .o1(m411));
 m_12 inst_452(.i1(m546),
              .i2(m401),
              .i3(m1454),
              .o1(m400));
 m_8 inst_453(.i1(m546),
             .i2(m401),
             .o1(m402));
 m_8 inst_454(.i1(m403),
             .i2(m404),
             .o1(m401));
 m_8 inst_455(.i1(m560),
             .i2(m561),
             .o1(m403));
 m_5 inst_456(.i1(m404),
             .o1(m405));
 m_6 inst_457(.i1(m1309),
             .i2(m406),
             .o1(m404));
 m_14 inst_458(.i1(i4[21]),
              .i2(i1[1]),
              .i3(m1308),
              .o1(m406));
 m_12 inst_459(.i1(i3[1]),
              .i2(m408),
              .i3(m410),
              .o1(m407));
 m_5 inst_460(.i1(m409),
             .o1(m408));
 m_20 inst_461(.i1(m560),
              .i2(m561),
              .o1(m409));
 m_10 inst_462(.i1(i3[1]),
              .i2(m421),
              .o1(m410));
 m_13 inst_463(.i1(m412),
              .i2(m618),
              .i3(m411),
              .o1(m553));
 m_10 inst_464(.i1(m1454),
              .i2(m549),
              .o1(m412));
 m_19 inst_465(.i1(m399),
              .i2(m400),
              .i3(o19),
              .i4(m413),
              .o1(m414));
 m_2 inst_466(.i1(m415),
             .i2(m414),
             .i3(o18),
             .o1(o5[17]));
 m_2 inst_467(.i1(m416),
             .i2(m415),
             .i3(o18),
             .o1(o5[9]));
 m_10 inst_468(.i1(m620),
              .i2(m413),
              .o1(m416));
 m_8 inst_469(.i1(o18),
             .i2(m416),
             .o1(o5[1]));
 m_10 inst_470(.i1(m620),
              .i2(m439),
              .o1(m415));
 m_12 inst_471(.i1(m605),
              .i2(m414),
              .i3(m417),
              .o1(o5[25]));
 m_14 inst_472(.i1(o19),
              .i2(m439),
              .i3(m537),
              .o1(m417));
 m_6 inst_473(.i1(m418),
             .i2(m423),
             .o1(m398));
 m_8 inst_474(.i1(m611),
             .i2(m419),
             .o1(m418));
 m_5 inst_475(.i1(m420),
             .o1(m419));
 m_6 inst_476(.i1(m611),
             .i2(m420),
             .o1(m421));
 m_6 inst_477(.i1(m1309),
             .i2(m422),
             .o1(m420));
 m_14 inst_478(.i1(i4[16]),
              .i2(i1[1]),
              .i3(m1308),
              .o1(m422));
 m_5 inst_479(.i1(m423),
             .o1(m424));
 m_18 inst_480(.i1(m611),
              .i2(m419),
              .i3(m424),
              .o1(m556));
 m_6 inst_481(.i1(m1309),
             .i2(m425),
             .o1(m423));
 m_14 inst_482(.i1(i4[17]),
              .i2(i1[1]),
              .i3(m1308),
              .o1(m425));
 m_12 inst_483(.i1(m397),
              .i2(m428),
              .i3(m620),
              .o1(m426));
 m_2 inst_484(.i1(m426),
             .i2(m504),
             .i3(o18),
             .o1(o5[21]));
 m_2 inst_485(.i1(m427),
             .i2(m426),
             .i3(o18),
             .o1(o5[13]));
 m_10 inst_486(.i1(m620),
              .i2(m522),
              .o1(m427));
 m_8 inst_487(.i1(o18),
             .i2(m427),
             .o1(o5[5]));
 m_8 inst_488(.i1(m1454),
             .i2(m429),
             .o1(m428));
 m_2 inst_489(.i1(m429),
             .i2(m430),
             .i3(m1454),
             .o1(m439));
 m_2 inst_490(.i1(m430),
             .i2(m431),
             .i3(m1454),
             .o1(m522));
 m_12 inst_491(.i1(i3[1]),
              .i2(m431),
              .i3(m432),
              .o1(m413));
 m_13 inst_492(.i1(i3[1]),
              .i2(m433),
              .i3(m434),
              .o1(m432));
 m_13 inst_493(.i1(i4[0]),
              .i2(i4[1]),
              .i3(m1309),
              .o1(m433));
 m_12 inst_494(.i1(m879),
              .i2(m232),
              .i3(m865),
              .o1(m434));
 m_6 inst_495(.i1(i4[5]),
             .i2(m435),
             .o1(m431));
 m_8 inst_496(.i1(m393),
             .i2(m232),
             .o1(m435));
 m_20 inst_497(.i1(m436),
              .i2(m437),
              .o1(m430));
 m_8 inst_498(.i1(m384),
             .i2(m385),
             .o1(m436));
 m_18 inst_499(.i1(m384),
              .i2(m385),
              .i3(m437),
              .o1(m348));
 m_6 inst_500(.i1(m614),
             .i2(m438),
             .o1(m437));
 m_8 inst_501(.i1(i4[9]),
             .i2(m1261),
             .o1(m438));
 m_20 inst_502(.i1(m440),
              .i2(m441),
              .o1(m429));
 m_8 inst_503(.i1(m513),
             .i2(m514),
             .o1(m440));
 m_18 inst_504(.i1(m513),
              .i2(m514),
              .i3(m441),
              .o1(m608));
 m_6 inst_505(.i1(m614),
             .i2(m442),
             .o1(m441));
 m_8 inst_506(.i1(i4[13]),
             .i2(m1261),
             .o1(m442));
 m_12 inst_507(.i1(m620),
              .i2(m396),
              .i3(m443),
              .o1(m478));
 m_13 inst_508(.i1(m444),
              .i2(m445),
              .i3(m443),
              .o1(m453));
 m_16 inst_509(.i1(i3[1]),
              .i2(m574),
              .o1(m444));
 m_10 inst_510(.i1(i3[1]),
              .i2(m446),
              .o1(m445));
 m_10 inst_511(.i1(m1454),
              .i2(m446),
              .o1(m447));
 m_12 inst_512(.i1(m1454),
              .i2(m543),
              .i3(m447),
              .o1(m455));
 m_8 inst_513(.i1(m474),
             .i2(m448),
             .o1(m446));
 m_5 inst_514(.i1(m449),
             .o1(m448));
 m_2 inst_515(.i1(m232),
             .i2(m1305),
             .i3(m450),
             .o1(m449));
 m_12 inst_516(.i1(i4[30]),
              .i2(m1302),
              .i3(m451),
              .o1(m450));
 m_13 inst_517(.i1(i4[7]),
              .i2(m1307),
              .i3(m451),
              .o1(m452));
 m_13 inst_518(.i1(m829),
              .i2(m1302),
              .i3(i1[0]),
              .o1(m451));
 m_12 inst_519(.i1(i3[1]),
              .i2(m574),
              .i3(m445),
              .o1(m528));
 m_8 inst_520(.i1(m454),
             .i2(m453),
             .o1(m456));
 m_16 inst_521(.i1(m537),
              .i2(m455),
              .o1(m454));
 m_13 inst_522(.i1(m456),
              .i2(m334),
              .i3(m603),
              .o1(m620));
 m_12 inst_523(.i1(m1454),
              .i2(m457),
              .i3(m477),
              .o1(m443));
 m_10 inst_524(.i1(m1454),
              .i2(m457),
              .o1(m458));
 m_12 inst_525(.i1(m1454),
              .i2(m459),
              .i3(m458),
              .o1(m537));
 m_6 inst_526(.i1(m460),
             .i2(m461),
             .o1(m459));
 m_10 inst_527(.i1(m460),
              .i2(m461),
              .o1(m336));
 m_6 inst_528(.i1(m1309),
             .i2(m462),
             .o1(m461));
 m_14 inst_529(.i1(i4[25]),
              .i2(i1[1]),
              .i3(m1308),
              .o1(m462));
 m_20 inst_530(.i1(m463),
              .i2(m475),
              .o1(m457));
 m_10 inst_531(.i1(m464),
              .i2(m471),
              .o1(m463));
 m_15 inst_532(.i1(m465),
              .i2(m466),
              .o1(m464));
 m_8 inst_533(.i1(m336),
             .i2(m337),
             .o1(m465));
 m_5 inst_534(.i1(m467),
             .o1(m466));
 m_12 inst_535(.i1(i4[31]),
              .i2(m468),
              .i3(m469),
              .o1(m467));
 m_10 inst_536(.i1(m659),
              .i2(i1[1]),
              .o1(m468));
 m_14 inst_537(.i1(i4[27]),
              .i2(i4[31]),
              .i3(m1302),
              .o1(m469));
 m_6 inst_538(.i1(m464),
             .i2(m471),
             .o1(m470));
 m_5 inst_539(.i1(m472),
             .o1(m471));
 m_12 inst_540(.i1(i4[31]),
              .i2(m666),
              .i3(m473),
              .o1(m472));
 m_14 inst_541(.i1(i4[28]),
              .i2(i4[31]),
              .i3(m1302),
              .o1(m473));
 m_16 inst_542(.i1(m463),
              .i2(m475),
              .o1(m474));
 m_12 inst_543(.i1(i4[29]),
              .i2(m1307),
              .i3(m476),
              .o1(m475));
 m_14 inst_544(.i1(i4[29]),
              .i2(i4[31]),
              .i3(m1302),
              .o1(m476));
 m_10 inst_545(.i1(m1454),
              .i2(m575),
              .o1(m477));
 m_8 inst_546(.i1(m479),
             .i2(m478),
             .o1(m496));
 m_5 inst_547(.i1(m479),
             .o1(m480));
 m_12 inst_548(.i1(m605),
              .i2(m481),
              .i3(m480),
              .o1(o5[24]));
 m_14 inst_549(.i1(o19),
              .i2(m378),
              .i3(m407),
              .o1(m481));
 m_2 inst_550(.i1(m482),
             .i2(m481),
             .i3(o18),
             .o1(o5[16]));
 m_2 inst_551(.i1(m483),
             .i2(m482),
             .i3(o18),
             .o1(o5[8]));
 m_8 inst_552(.i1(o18),
             .i2(m483),
             .o1(o5[0]));
 m_12 inst_553(.i1(m620),
              .i2(m484),
              .i3(m485),
              .o1(m479));
 m_5 inst_554(.i1(m381),
             .o1(m484));
 m_13 inst_555(.i1(m486),
              .i2(m485),
              .i3(m487),
              .o1(m602));
 m_5 inst_556(.i1(m531),
             .o1(m486));
 m_8 inst_557(.i1(m544),
             .i2(m488),
             .o1(m487));
 m_12 inst_558(.i1(m1454),
              .i2(m489),
              .i3(m495),
              .o1(m485));
 m_10 inst_559(.i1(m1454),
              .i2(m489),
              .o1(m490));
 m_12 inst_560(.i1(m1454),
              .i2(m408),
              .i3(m490),
              .o1(m506));
 m_20 inst_561(.i1(m491),
              .i2(m492),
              .o1(m489));
 m_8 inst_562(.i1(m491),
             .i2(m492),
             .o1(m460));
 m_12 inst_563(.i1(i4[31]),
              .i2(m493),
              .i3(m494),
              .o1(m492));
 m_10 inst_564(.i1(m703),
              .i2(i1[1]),
              .o1(m493));
 m_14 inst_565(.i1(i4[24]),
              .i2(i4[31]),
              .i3(m1302),
              .o1(m494));
 m_10 inst_566(.i1(m1454),
              .i2(m470),
              .o1(m495));
 m_13 inst_567(.i1(m497),
              .i2(m604),
              .i3(m496),
              .o1(m502));
 m_14 inst_568(.i1(o19),
              .i2(m518),
              .i3(m455),
              .o1(m497));
 m_12 inst_569(.i1(m605),
              .i2(m498),
              .i3(m497),
              .o1(o5[27]));
 m_2 inst_570(.i1(m499),
             .i2(m498),
             .i3(o18),
             .o1(o5[19]));
 m_2 inst_571(.i1(m500),
             .i2(m499),
             .i3(o18),
             .o1(o5[11]));
 m_8 inst_572(.i1(o18),
             .i2(m500),
             .o1(o5[3]));
 m_16 inst_573(.i1(m478),
              .i2(m501),
              .o1(o5[29]));
 m_18 inst_574(.i1(m502),
              .i2(m503),
              .i3(m504),
              .o1(m501));
 m_16 inst_575(.i1(m502),
              .i2(m503),
              .o1(m605));
 m_14 inst_576(.i1(o19),
              .i2(m522),
              .i3(m505),
              .o1(m504));
 m_18 inst_577(.i1(m505),
              .i2(m506),
              .i3(m554),
              .o1(m507));
 m_13 inst_578(.i1(m624),
              .i2(m625),
              .i3(m507),
              .o1(m488));
 m_12 inst_579(.i1(i3[1]),
              .i2(m459),
              .i3(m508),
              .o1(m505));
 m_10 inst_580(.i1(i3[1]),
              .i2(m402),
              .o1(m508));
 m_5 inst_581(.i1(m510),
             .o1(m509));
 m_10 inst_582(.i1(m620),
              .i2(m510),
              .o1(m511));
 m_2 inst_583(.i1(m388),
             .i2(m511),
             .i3(o18),
             .o1(o5[12]));
 m_12 inst_584(.i1(m1454),
              .i2(m512),
              .i3(m516),
              .o1(m510));
 m_6 inst_585(.i1(m513),
             .i2(m514),
             .o1(m512));
 m_6 inst_586(.i1(m614),
             .i2(m515),
             .o1(m514));
 m_8 inst_587(.i1(i4[12]),
             .i2(m1261),
             .o1(m515));
 m_10 inst_588(.i1(m1454),
              .i2(m421),
              .o1(m516));
 m_8 inst_589(.i1(m518),
             .i2(m519),
             .o1(m517));
 m_10 inst_590(.i1(m620),
              .i2(m518),
              .o1(m499));
 m_13 inst_591(.i1(m520),
              .i2(m521),
              .i3(m525),
              .o1(m519));
 m_5 inst_592(.i1(m627),
             .o1(m520));
 m_8 inst_593(.i1(m522),
             .i2(m523),
             .o1(m521));
 m_12 inst_594(.i1(i3[1]),
              .i2(m1323),
              .i3(m524),
              .o1(m523));
 m_8 inst_595(.i1(m1322),
             .i2(m413),
             .o1(m524));
 m_8 inst_596(.i1(m439),
             .i2(m357),
             .o1(m525));
 m_8 inst_597(.i1(m527),
             .i2(m569),
             .o1(m526));
 m_14 inst_598(.i1(o19),
              .i2(m527),
              .i3(m528),
              .o1(m529));
 m_13 inst_599(.i1(m529),
              .i2(m530),
              .i3(m533),
              .o1(m503));
 m_14 inst_600(.i1(o19),
              .i2(m510),
              .i3(m531),
              .o1(m530));
 m_2 inst_601(.i1(m470),
             .i2(m576),
             .i3(i3[1]),
             .o1(m531));
 m_12 inst_602(.i1(m605),
              .i2(m532),
              .i3(m530),
              .o1(o5[28]));
 m_14 inst_603(.i1(o19),
              .i2(m387),
              .i3(m506),
              .o1(m532));
 m_2 inst_604(.i1(m511),
             .i2(m532),
             .i3(o18),
             .o1(o5[20]));
 m_8 inst_605(.i1(m339),
             .i2(m534),
             .o1(m533));
 m_12 inst_606(.i1(m620),
              .i2(m535),
              .i3(m536),
              .o1(m534));
 m_5 inst_607(.i1(m439),
             .o1(m535));
 m_5 inst_608(.i1(m537),
             .o1(m536));
 m_12 inst_609(.i1(m605),
              .i2(m539),
              .i3(m529),
              .o1(o5[31]));
 m_10 inst_610(.i1(m620),
              .i2(m527),
              .o1(m538));
 m_2 inst_611(.i1(m538),
             .i2(m539),
             .i3(o18),
             .o1(o5[23]));
 m_14 inst_612(.i1(o19),
              .i2(m359),
              .i3(m544),
              .o1(m539));
 m_2 inst_613(.i1(m540),
             .i2(m538),
             .i3(o18),
             .o1(o5[15]));
 m_10 inst_614(.i1(m620),
              .i2(m359),
              .o1(m540));
 m_8 inst_615(.i1(o18),
             .i2(m540),
             .o1(o5[7]));
 m_12 inst_616(.i1(i3[1]),
              .i2(m541),
              .i3(m564),
              .o1(m527));
 m_2 inst_617(.i1(m542),
             .i2(m541),
             .i3(m1454),
             .o1(m552));
 m_2 inst_618(.i1(m543),
             .i2(m542),
             .i3(m1454),
             .o1(m544));
 m_6 inst_619(.i1(m465),
             .i2(m466),
             .o1(m543));
 m_6 inst_620(.i1(m545),
             .i2(m550),
             .o1(m542));
 m_15 inst_621(.i1(m546),
              .i2(m547),
              .o1(m545));
 m_8 inst_622(.i1(m545),
             .i2(m548),
             .o1(m549));
 m_8 inst_623(.i1(m546),
             .i2(m547),
             .o1(m548));
 m_10 inst_624(.i1(i3[1]),
              .i2(m549),
              .o1(m625));
 m_13 inst_625(.i1(m546),
              .i2(m547),
              .i3(m550),
              .o1(m491));
 m_6 inst_626(.i1(m1309),
             .i2(m551),
             .o1(m550));
 m_14 inst_627(.i1(i4[23]),
              .i2(i1[1]),
              .i3(m1308),
              .o1(m551));
 m_14 inst_628(.i1(o19),
              .i2(m379),
              .i3(m552),
              .o1(m498));
 m_16 inst_629(.i1(m552),
              .i2(m553),
              .o1(m554));
 m_6 inst_630(.i1(m555),
             .i2(m559),
             .o1(m541));
 m_15 inst_631(.i1(m556),
              .i2(m557),
              .o1(m555));
 m_14 inst_632(.i1(i4[18]),
              .i2(i4[31]),
              .i3(m558),
              .o1(m557));
 m_12 inst_633(.i1(i4[18]),
              .i2(i4[31]),
              .i3(i1[1]),
              .o1(m558));
 m_13 inst_634(.i1(m556),
              .i2(m557),
              .i3(m559),
              .o1(m560));
 m_18 inst_635(.i1(m560),
              .i2(m561),
              .i3(m405),
              .o1(m546));
 m_12 inst_636(.i1(i4[20]),
              .i2(i4[31]),
              .i3(m562),
              .o1(m561));
 m_14 inst_637(.i1(i4[20]),
              .i2(i4[31]),
              .i3(m1302),
              .o1(m562));
 m_6 inst_638(.i1(m1309),
             .i2(m563),
             .o1(m559));
 m_14 inst_639(.i1(i4[19]),
              .i2(i1[1]),
              .i3(m1308),
              .o1(m563));
 m_10 inst_640(.i1(i3[1]),
              .i2(m565),
              .o1(m564));
 m_10 inst_641(.i1(m1454),
              .i2(m565),
              .o1(m566));
 m_12 inst_642(.i1(m1454),
              .i2(m360),
              .i3(m566),
              .o1(m518));
 m_8 inst_643(.i1(m567),
             .i2(m568),
             .o1(m565));
 m_5 inst_644(.i1(m611),
             .o1(m567));
 m_14 inst_645(.i1(m608),
              .i2(m612),
              .i3(m609),
              .o1(m568));
 m_14 inst_646(.i1(o19),
              .i2(m569),
              .i3(m570),
              .o1(m604));
 m_2 inst_647(.i1(m571),
             .i2(m573),
             .i3(i3[1]),
             .o1(m570));
 m_10 inst_648(.i1(m1454),
              .i2(m571),
              .o1(m572));
 m_6 inst_649(.i1(m474),
             .i2(m448),
             .o1(m571));
 m_2 inst_650(.i1(m573),
             .i2(m574),
             .i3(m1459),
             .o1(o4[24]));
 m_2 inst_651(.i1(i10[26]),
             .i2(i11[26]),
             .i3(m1203),
             .o1(m574));
 m_2 inst_652(.i1(m575),
             .i2(m573),
             .i3(m1459),
             .o1(o4[23]));
 m_2 inst_653(.i1(m576),
             .i2(m575),
             .i3(m1459),
             .o1(o4[22]));
 m_2 inst_654(.i1(m577),
             .i2(m576),
             .i3(m1459),
             .o1(o4[21]));
 m_2 inst_655(.i1(m578),
             .i2(m577),
             .i3(m1459),
             .o1(o4[20]));
 m_2 inst_656(.i1(m579),
             .i2(m578),
             .i3(m1459),
             .o1(o4[19]));
 m_2 inst_657(.i1(m580),
             .i2(m579),
             .i3(m1459),
             .o1(o4[18]));
 m_2 inst_658(.i1(m581),
             .i2(m580),
             .i3(m1459),
             .o1(o4[17]));
 m_2 inst_659(.i1(m582),
             .i2(m581),
             .i3(m1459),
             .o1(o4[16]));
 m_2 inst_660(.i1(m583),
             .i2(m582),
             .i3(m1459),
             .o1(o4[15]));
 m_2 inst_661(.i1(m584),
             .i2(m583),
             .i3(m1459),
             .o1(o4[14]));
 m_2 inst_662(.i1(m585),
             .i2(m584),
             .i3(m1459),
             .o1(o4[13]));
 m_2 inst_663(.i1(m586),
             .i2(m585),
             .i3(m1459),
             .o1(o4[12]));
 m_2 inst_664(.i1(m587),
             .i2(m586),
             .i3(m1459),
             .o1(o4[11]));
 m_2 inst_665(.i1(m588),
             .i2(m587),
             .i3(m1459),
             .o1(o4[10]));
 m_2 inst_666(.i1(m589),
             .i2(m588),
             .i3(m1459),
             .o1(o4[9]));
 m_2 inst_667(.i1(m590),
             .i2(m589),
             .i3(m1459),
             .o1(o4[8]));
 m_2 inst_668(.i1(m591),
             .i2(m590),
             .i3(m1459),
             .o1(o4[7]));
 m_2 inst_669(.i1(m592),
             .i2(m591),
             .i3(m1459),
             .o1(o4[6]));
 m_2 inst_670(.i1(m593),
             .i2(m592),
             .i3(m1459),
             .o1(o4[5]));
 m_2 inst_671(.i1(m594),
             .i2(m593),
             .i3(m1459),
             .o1(o4[4]));
 m_2 inst_672(.i1(m595),
             .i2(m594),
             .i3(m1459),
             .o1(o4[3]));
 m_2 inst_673(.i1(m596),
             .i2(m595),
             .i3(m1459),
             .o1(o4[2]));
 m_2 inst_674(.i1(m597),
             .i2(m596),
             .i3(m1459),
             .o1(o4[1]));
 m_2 inst_675(.i1(i10[2]),
             .i2(i11[2]),
             .i3(m1203),
             .o1(m597));
 m_12 inst_676(.i1(m597),
              .i2(m1459),
              .i3(m598),
              .o1(o4[0]));
 m_12 inst_677(.i1(i11[0]),
              .i2(m599),
              .i3(m600),
              .o1(m598));
 m_16 inst_678(.i1(i11[1]),
              .i2(m1203),
              .o1(m599));
 m_10 inst_679(.i1(m1203),
              .i2(m601),
              .o1(m600));
 m_8 inst_680(.i1(i10[0]),
             .i2(i10[1]),
             .o1(m601));
 m_2 inst_681(.i1(i10[3]),
             .i2(i11[3]),
             .i3(m1203),
             .o1(m596));
 m_2 inst_682(.i1(i10[4]),
             .i2(i11[4]),
             .i3(m1203),
             .o1(m595));
 m_2 inst_683(.i1(i10[5]),
             .i2(i11[5]),
             .i3(m1203),
             .o1(m594));
 m_2 inst_684(.i1(i10[6]),
             .i2(i11[6]),
             .i3(m1203),
             .o1(m593));
 m_2 inst_685(.i1(i10[7]),
             .i2(i11[7]),
             .i3(m1203),
             .o1(m592));
 m_2 inst_686(.i1(i10[8]),
             .i2(i11[8]),
             .i3(m1203),
             .o1(m591));
 m_2 inst_687(.i1(i10[9]),
             .i2(i11[9]),
             .i3(m1203),
             .o1(m590));
 m_2 inst_688(.i1(i10[10]),
             .i2(i11[10]),
             .i3(m1203),
             .o1(m589));
 m_2 inst_689(.i1(i10[11]),
             .i2(i11[11]),
             .i3(m1203),
             .o1(m588));
 m_2 inst_690(.i1(i10[12]),
             .i2(i11[12]),
             .i3(m1203),
             .o1(m587));
 m_2 inst_691(.i1(i10[13]),
             .i2(i11[13]),
             .i3(m1203),
             .o1(m586));
 m_2 inst_692(.i1(i10[14]),
             .i2(i11[14]),
             .i3(m1203),
             .o1(m585));
 m_2 inst_693(.i1(i10[15]),
             .i2(i11[15]),
             .i3(m1203),
             .o1(m584));
 m_2 inst_694(.i1(i10[16]),
             .i2(i11[16]),
             .i3(m1203),
             .o1(m583));
 m_2 inst_695(.i1(i10[17]),
             .i2(i11[17]),
             .i3(m1203),
             .o1(m582));
 m_2 inst_696(.i1(i10[18]),
             .i2(i11[18]),
             .i3(m1203),
             .o1(m581));
 m_2 inst_697(.i1(i10[19]),
             .i2(i11[19]),
             .i3(m1203),
             .o1(m580));
 m_2 inst_698(.i1(i10[20]),
             .i2(i11[20]),
             .i3(m1203),
             .o1(m579));
 m_2 inst_699(.i1(i10[21]),
             .i2(i11[21]),
             .i3(m1203),
             .o1(m578));
 m_2 inst_700(.i1(i10[22]),
             .i2(i11[22]),
             .i3(m1203),
             .o1(m577));
 m_2 inst_701(.i1(i10[23]),
             .i2(i11[23]),
             .i3(m1203),
             .o1(m576));
 m_2 inst_702(.i1(i10[24]),
             .i2(i11[24]),
             .i3(m1203),
             .o1(m575));
 m_2 inst_703(.i1(i10[25]),
             .i2(i11[25]),
             .i3(m1203),
             .o1(m573));
 m_8 inst_704(.i1(m570),
             .i2(m602),
             .o1(m603));
 m_12 inst_705(.i1(m605),
              .i2(m622),
              .i3(m604),
              .o1(o5[30]));
 m_5 inst_706(.i1(m605),
             .o1(o18));
 m_14 inst_707(.i1(i3[1]),
              .i2(m606),
              .i3(m616),
              .o1(m569));
 m_10 inst_708(.i1(m1454),
              .i2(m606),
              .o1(m607));
 m_6 inst_709(.i1(m608),
             .i2(m612),
             .o1(m606));
 m_13 inst_710(.i1(m608),
              .i2(m612),
              .i3(m609),
              .o1(m611));
 m_6 inst_711(.i1(m614),
             .i2(m610),
             .o1(m609));
 m_12 inst_712(.i1(i1[1]),
              .i2(i1[0]),
              .i3(m829),
              .o1(m610));
 m_5 inst_713(.i1(m613),
             .o1(m612));
 m_6 inst_714(.i1(m614),
             .i2(m615),
             .o1(m613));
 m_8 inst_715(.i1(i4[14]),
             .i2(m1261),
             .o1(m615));
 m_8 inst_716(.i1(i3[1]),
             .i2(m617),
             .o1(m616));
 m_10 inst_717(.i1(i3[1]),
              .i2(m617),
              .o1(m618));
 m_10 inst_718(.i1(m412),
              .i2(m618),
              .o1(m355));
 m_8 inst_719(.i1(m555),
             .i2(m619),
             .o1(m617));
 m_8 inst_720(.i1(m556),
             .i2(m557),
             .o1(m619));
 m_10 inst_721(.i1(m620),
              .i2(m569),
              .o1(m621));
 m_2 inst_722(.i1(m621),
             .i2(m622),
             .i3(o18),
             .o1(o5[22]));
 m_14 inst_723(.i1(o19),
              .i2(m627),
              .i3(m623),
              .o1(m622));
 m_10 inst_724(.i1(m624),
              .i2(m625),
              .o1(m623));
 m_2 inst_725(.i1(m626),
             .i2(m621),
             .i3(o18),
             .o1(o5[14]));
 m_10 inst_726(.i1(m620),
              .i2(m627),
              .o1(m626));
 m_8 inst_727(.i1(o18),
             .i2(m626),
             .o1(o5[6]));
 m_12 inst_728(.i1(m628),
              .i2(m747),
              .i3(m326),
              .o1(o15));
 m_13 inst_729(.i1(m629),
              .i2(m673),
              .i3(m746),
              .o1(m628));
 m_8 inst_730(.i1(m630),
             .i2(m631),
             .o1(m629));
 m_8 inst_731(.i1(m631),
             .i2(m311),
             .o1(m632));
 m_12 inst_732(.i1(m632),
              .i2(m633),
              .i3(m635),
              .o1(m637));
 m_19 inst_733(.i1(m301),
              .i2(m311),
              .i3(m634),
              .i4(m646),
              .o1(m633));
 m_6 inst_734(.i1(m636),
             .i2(m746),
             .o1(m635));
 m_18 inst_735(.i1(m1195),
              .i2(m1196),
              .i3(m637),
              .o1(m281));
 m_8 inst_736(.i1(m638),
             .i2(i5[29]),
             .o1(m631));
 m_5 inst_737(.i1(i4[29]),
             .o1(m638));
 m_10 inst_738(.i1(m638),
              .i2(i5[29]),
              .o1(m301));
 m_12 inst_739(.i1(m638),
              .i2(i5[29]),
              .i3(m303),
              .o1(m639));
 m_14 inst_740(.i1(m639),
              .i2(m672),
              .i3(m640),
              .o1(m641));
 m_20 inst_741(.i1(m636),
              .i2(m746),
              .o1(m640));
 m_13 inst_742(.i1(m642),
              .i2(m643),
              .i3(m641),
              .o1(m295));
 m_14 inst_743(.i1(m642),
              .i2(m643),
              .i3(i3[1]),
              .o1(m240));
 m_5 inst_744(.i1(m642),
             .o1(m1195));
 m_10 inst_745(.i1(m931),
              .i2(i5[30]),
              .o1(m642));
 m_12 inst_746(.i1(i4[30]),
              .i2(m644),
              .i3(m643),
              .o1(m1198));
 m_19 inst_747(.i1(i4[30]),
              .i2(m644),
              .i3(m301),
              .i4(m302),
              .o1(m1196));
 m_5 inst_748(.i1(i5[30]),
             .o1(m644));
 m_10 inst_749(.i1(m931),
              .i2(m644),
              .o1(o17[30]));
 m_17 inst_750(.i1(m931),
              .i2(i5[30]),
              .i3(m630),
              .i4(m310),
              .o1(m643));
 m_16 inst_751(.i1(m630),
              .i2(m631),
              .o1(m645));
 m_14 inst_752(.i1(m646),
              .i2(m647),
              .i3(m645),
              .o1(m310));
 m_10 inst_753(.i1(m665),
              .i2(i5[28]),
              .o1(m646));
 m_12 inst_754(.i1(m656),
              .i2(m648),
              .i3(m649),
              .o1(m647));
 m_14 inst_755(.i1(m740),
              .i2(m663),
              .i3(m658),
              .o1(m648));
 m_10 inst_756(.i1(i4[28]),
              .i2(m650),
              .o1(m649));
 m_5 inst_757(.i1(i5[28]),
             .o1(m650));
 m_8 inst_758(.i1(i4[28]),
             .i2(m650),
             .o1(m653));
 m_12 inst_759(.i1(m1195),
              .i2(m1196),
              .i3(m650),
              .o1(m651));
 m_12 inst_760(.i1(i4[28]),
              .i2(m1198),
              .i3(m651),
              .o1(m652));
 m_5 inst_761(.i1(m652),
             .o1(o17[28]));
 m_18 inst_762(.i1(m629),
              .i2(m653),
              .i3(m654),
              .o1(m316));
 m_14 inst_763(.i1(m655),
              .i2(m661),
              .i3(m664),
              .o1(m654));
 m_5 inst_764(.i1(m655),
             .o1(m656));
 m_10 inst_765(.i1(m655),
              .i2(m657),
              .o1(m658));
 m_5 inst_766(.i1(m658),
             .o1(m739));
 m_10 inst_767(.i1(m659),
              .i2(i5[27]),
              .o1(m655));
 m_5 inst_768(.i1(i4[27]),
             .o1(m659));
 m_12 inst_769(.i1(m659),
              .i2(m1198),
              .i3(m660),
              .o1(o17[27]));
 m_12 inst_770(.i1(m1195),
              .i2(m1196),
              .i3(i5[27]),
              .o1(m660));
 m_15 inst_771(.i1(m661),
              .i2(m662),
              .o1(m239));
 m_13 inst_772(.i1(m658),
              .i2(m740),
              .i3(m663),
              .o1(m662));
 m_8 inst_773(.i1(m664),
             .i2(m653),
             .o1(m746));
 m_8 inst_774(.i1(m665),
             .i2(i5[28]),
             .o1(m664));
 m_5 inst_775(.i1(i4[28]),
             .o1(m665));
 m_10 inst_776(.i1(m665),
              .i2(i1[1]),
              .o1(m666));
 m_18 inst_777(.i1(m664),
              .i2(m667),
              .i3(m668),
              .o1(m671));
 m_5 inst_778(.i1(m657),
             .o1(m667));
 m_14 inst_779(.i1(m713),
              .i2(m669),
              .i3(m658),
              .o1(m668));
 m_12 inst_780(.i1(m670),
              .i2(m710),
              .i3(m740),
              .o1(m669));
 m_8 inst_781(.i1(m742),
             .i2(i5[25]),
             .o1(m670));
 m_17 inst_782(.i1(m630),
              .i2(m303),
              .i3(m671),
              .i4(m653),
              .o1(m672));
 m_12 inst_783(.i1(m653),
              .i2(m654),
              .i3(m629),
              .o1(m302));
 m_12 inst_784(.i1(m702),
              .i2(m704),
              .i3(m673),
              .o1(m707));
 m_12 inst_785(.i1(m674),
              .i2(m688),
              .i3(m673),
              .o1(m692));
 m_8 inst_786(.i1(i4[24]),
             .i2(m675),
             .o1(m674));
 m_5 inst_787(.i1(i5[24]),
             .o1(m675));
 m_12 inst_788(.i1(m1195),
              .i2(m1196),
              .i3(m675),
              .o1(m676));
 m_12 inst_789(.i1(i4[24]),
              .i2(m1198),
              .i3(m676),
              .o1(m677));
 m_5 inst_790(.i1(m677),
             .o1(o17[24]));
 m_10 inst_791(.i1(m691),
              .i2(m677),
              .o1(m678));
 m_12 inst_792(.i1(o17[25]),
              .i2(m678),
              .i3(o17[26]),
              .o1(m679));
 m_15 inst_793(.i1(m679),
              .i2(m718),
              .o1(m680));
 m_12 inst_794(.i1(m685),
              .i2(m680),
              .i3(m681),
              .o1(o6[28]));
 m_12 inst_795(.i1(i18[26]),
              .i2(o13),
              .i3(i18[30]),
              .o1(m681));
 m_20 inst_796(.i1(o17[25]),
              .i2(m678),
              .o1(m682));
 m_12 inst_797(.i1(m685),
              .i2(m682),
              .i3(m683),
              .o1(o6[27]));
 m_12 inst_798(.i1(i18[26]),
              .i2(o13),
              .i3(i18[29]),
              .o1(m683));
 m_20 inst_799(.i1(m691),
              .i2(m677),
              .o1(m684));
 m_12 inst_800(.i1(m685),
              .i2(m684),
              .i3(m687),
              .o1(o6[26]));
 m_12 inst_801(.i1(o17[23]),
              .i2(m685),
              .i3(m686),
              .o1(o6[25]));
 m_12 inst_802(.i1(i18[26]),
              .i2(o13),
              .i3(i18[27]),
              .o1(m686));
 m_16 inst_803(.i1(i18[26]),
              .i2(o13),
              .o1(m685));
 m_12 inst_804(.i1(i18[26]),
              .i2(o13),
              .i3(i18[28]),
              .o1(m687));
 m_14 inst_805(.i1(i4[23]),
              .i2(m689),
              .i3(m706),
              .o1(m688));
 m_5 inst_806(.i1(i5[23]),
             .o1(m689));
 m_8 inst_807(.i1(i4[23]),
             .i2(m689),
             .o1(m183));
 m_12 inst_808(.i1(m1195),
              .i2(m1196),
              .i3(m689),
              .o1(m690));
 m_12 inst_809(.i1(i4[23]),
              .i2(m1198),
              .i3(m690),
              .o1(m691));
 m_5 inst_810(.i1(m691),
             .o1(o17[23]));
 m_6 inst_811(.i1(i18[27]),
             .i2(m691),
             .o1(m1326));
 m_20 inst_812(.i1(i18[27]),
              .i2(m691),
              .o1(m1424));
 m_14 inst_813(.i1(m693),
              .i2(m692),
              .i3(m695),
              .o1(m699));
 m_5 inst_814(.i1(m694),
             .o1(m693));
 m_8 inst_815(.i1(i4[25]),
             .i2(m700),
             .o1(m694));
 m_12 inst_816(.i1(m694),
              .i2(m293),
              .i3(m713),
              .o1(m663));
 m_8 inst_817(.i1(m695),
             .i2(m696),
             .o1(m877));
 m_8 inst_818(.i1(i4[26]),
             .i2(m714),
             .o1(m696));
 m_8 inst_819(.i1(m697),
             .i2(i5[26]),
             .o1(m695));
 m_5 inst_820(.i1(i4[26]),
             .o1(m697));
 m_10 inst_821(.i1(m697),
              .i2(i1[1]),
              .o1(m698));
 m_10 inst_822(.i1(m697),
              .i2(i5[26]),
              .o1(m740));
 m_12 inst_823(.i1(m696),
              .i2(m699),
              .i3(m739),
              .o1(m661));
 m_12 inst_824(.i1(i4[25]),
              .i2(m700),
              .i3(m692),
              .o1(m701));
 m_5 inst_825(.i1(i5[25]),
             .o1(m700));
 m_20 inst_826(.i1(m701),
              .i2(m877),
              .o1(m237));
 m_8 inst_827(.i1(m703),
             .i2(i5[24]),
             .o1(m702));
 m_5 inst_828(.i1(i4[24]),
             .o1(m703));
 m_14 inst_829(.i1(m705),
              .i2(i5[23]),
              .i3(m706),
              .o1(m704));
 m_5 inst_830(.i1(i4[23]),
             .o1(m705));
 m_8 inst_831(.i1(m705),
             .i2(i5[23]),
             .o1(m182));
 m_20 inst_832(.i1(i4[24]),
              .i2(i5[24]),
              .o1(m706));
 m_15 inst_833(.i1(m707),
              .i2(m708),
              .o1(m712));
 m_13 inst_834(.i1(m291),
              .i2(m709),
              .i3(m711),
              .o1(m708));
 m_14 inst_835(.i1(m709),
              .i2(m711),
              .i3(m291),
              .o1(m710));
 m_10 inst_836(.i1(i4[24]),
              .i2(m675),
              .o1(m709));
 m_12 inst_837(.i1(i4[23]),
              .i2(m689),
              .i3(m288),
              .o1(m711));
 m_13 inst_838(.i1(m713),
              .i2(m734),
              .i3(m707),
              .o1(m735));
 m_10 inst_839(.i1(i4[26]),
              .i2(m714),
              .o1(m713));
 m_5 inst_840(.i1(i5[26]),
             .o1(m714));
 m_12 inst_841(.i1(m1195),
              .i2(m1196),
              .i3(m714),
              .o1(m715));
 m_12 inst_842(.i1(i4[26]),
              .i2(m1198),
              .i3(m715),
              .o1(m716));
 m_5 inst_843(.i1(m716),
             .o1(o17[26]));
 m_10 inst_844(.i1(m716),
              .i2(m717),
              .o1(m718));
 m_8 inst_845(.i1(o17[25]),
             .i2(m678),
             .o1(m717));
 m_8 inst_846(.i1(o17[27]),
             .i2(m718),
             .o1(m719));
 m_15 inst_847(.i1(m652),
              .i2(m719),
              .o1(m720));
 m_10 inst_848(.i1(m721),
              .i2(m720),
              .o1(m724));
 m_5 inst_849(.i1(m721),
             .o1(o17[29]));
 m_12 inst_850(.i1(i4[29]),
              .i2(m1198),
              .i3(m722),
              .o1(m721));
 m_12 inst_851(.i1(m1195),
              .i2(m1196),
              .i3(m723),
              .o1(m722));
 m_5 inst_852(.i1(i5[29]),
             .o1(m723));
 m_8 inst_853(.i1(i4[29]),
             .i2(m723),
             .o1(m630));
 m_20 inst_854(.i1(o17[30]),
              .i2(m724),
              .o1(m725));
 m_12 inst_855(.i1(m685),
              .i2(m725),
              .i3(m726),
              .o1(o6[32]));
 m_12 inst_856(.i1(i18[26]),
              .i2(o13),
              .i3(i18[34]),
              .o1(m726));
 m_6 inst_857(.i1(o17[29]),
             .i2(m720),
             .o1(m727));
 m_12 inst_858(.i1(m685),
              .i2(m727),
              .i3(m728),
              .o1(o6[31]));
 m_12 inst_859(.i1(i18[26]),
              .i2(o13),
              .i3(i18[33]),
              .o1(m728));
 m_8 inst_860(.i1(m652),
             .i2(m719),
             .o1(m729));
 m_8 inst_861(.i1(m729),
             .i2(m720),
             .o1(m730));
 m_12 inst_862(.i1(m685),
              .i2(m730),
              .i3(m731),
              .o1(o6[30]));
 m_12 inst_863(.i1(i18[26]),
              .i2(o13),
              .i3(i18[32]),
              .o1(m731));
 m_20 inst_864(.i1(o17[27]),
              .i2(m718),
              .o1(m732));
 m_12 inst_865(.i1(m685),
              .i2(m732),
              .i3(m733),
              .o1(o6[29]));
 m_12 inst_866(.i1(i18[26]),
              .i2(o13),
              .i3(i18[31]),
              .o1(m733));
 m_10 inst_867(.i1(i4[25]),
              .i2(m700),
              .o1(m734));
 m_14 inst_868(.i1(m740),
              .i2(m735),
              .i3(m739),
              .o1(m736));
 m_8 inst_869(.i1(m668),
             .i2(m736),
             .o1(m737));
 m_16 inst_870(.i1(i3[1]),
              .i2(m737),
              .o1(m738));
 m_12 inst_871(.i1(m295),
              .i2(m738),
              .i3(m284),
              .o1(m256));
 m_13 inst_872(.i1(m739),
              .i2(m740),
              .i3(m735),
              .o1(m741));
 m_13 inst_873(.i1(m649),
              .i2(m657),
              .i3(m741),
              .o1(m634));
 m_12 inst_874(.i1(m659),
              .i2(i5[27]),
              .i3(m741),
              .o1(m636));
 m_12 inst_875(.i1(m742),
              .i2(i5[25]),
              .i3(m707),
              .o1(m744));
 m_5 inst_876(.i1(i4[25]),
             .o1(m742));
 m_12 inst_877(.i1(m742),
              .i2(m1198),
              .i3(m743),
              .o1(o17[25]));
 m_12 inst_878(.i1(m1195),
              .i2(m1196),
              .i3(i5[25]),
              .o1(m743));
 m_20 inst_879(.i1(m744),
              .i2(m877),
              .o1(m745));
 m_6 inst_880(.i1(i4[25]),
             .i2(i5[25]),
             .o1(m673));
 m_13 inst_881(.i1(m748),
              .i2(m837),
              .i3(m881),
              .o1(m747));
 m_8 inst_882(.i1(m749),
             .i2(m779),
             .o1(m748));
 m_14 inst_883(.i1(m750),
              .i2(m751),
              .i3(m749),
              .o1(m754));
 m_13 inst_884(.i1(m780),
              .i2(m803),
              .i3(m793),
              .o1(m750));
 m_12 inst_885(.i1(m752),
              .i2(i5[11]),
              .i3(m781),
              .o1(m751));
 m_5 inst_886(.i1(i4[11]),
             .o1(m752));
 m_12 inst_887(.i1(m752),
              .i2(m185),
              .i3(m753),
              .o1(o20[12]));
 m_12 inst_888(.i1(m182),
              .i2(m183),
              .i3(i4[12]),
              .o1(m753));
 m_14 inst_889(.i1(m755),
              .i2(m774),
              .i3(m754),
              .o1(m832));
 m_10 inst_890(.i1(m755),
              .i2(m769),
              .o1(m749));
 m_8 inst_891(.i1(m756),
             .i2(m765),
             .o1(m755));
 m_17 inst_892(.i1(i4[14]),
              .i2(m757),
              .i3(i4[15]),
              .i4(m761),
              .o1(m756));
 m_5 inst_893(.i1(i5[14]),
             .o1(m757));
 m_12 inst_894(.i1(m757),
              .i2(m1200),
              .i3(m758),
              .o1(o21[14]));
 m_10 inst_895(.i1(i5[13]),
              .i2(m1200),
              .o1(m758));
 m_12 inst_896(.i1(m1195),
              .i2(m1196),
              .i3(m757),
              .o1(m759));
 m_12 inst_897(.i1(i4[14]),
              .i2(m1198),
              .i3(m759),
              .o1(m760));
 m_5 inst_898(.i1(m760),
             .o1(o17[14]));
 m_5 inst_899(.i1(i5[15]),
             .o1(m761));
 m_12 inst_900(.i1(m761),
              .i2(m1200),
              .i3(m762),
              .o1(o21[15]));
 m_10 inst_901(.i1(i5[14]),
              .i2(m1200),
              .o1(m762));
 m_12 inst_902(.i1(m1195),
              .i2(m1196),
              .i3(m761),
              .o1(m763));
 m_12 inst_903(.i1(i4[15]),
              .i2(m1198),
              .i3(m763),
              .o1(m764));
 m_5 inst_904(.i1(m764),
             .o1(o17[15]));
 m_12 inst_905(.i1(m766),
              .i2(i5[13]),
              .i3(m768),
              .o1(m765));
 m_5 inst_906(.i1(i4[13]),
             .o1(m766));
 m_12 inst_907(.i1(m766),
              .i2(m185),
              .i3(m767),
              .o1(o20[14]));
 m_12 inst_908(.i1(m182),
              .i2(m183),
              .i3(i4[14]),
              .o1(m767));
 m_19 inst_909(.i1(i4[14]),
              .i2(m757),
              .i3(i4[15]),
              .i4(m761),
              .o1(m768));
 m_14 inst_910(.i1(i4[12]),
              .i2(m770),
              .i3(m774),
              .o1(m769));
 m_5 inst_911(.i1(i5[12]),
             .o1(m770));
 m_12 inst_912(.i1(m770),
              .i2(m1200),
              .i3(m771),
              .o1(o21[12]));
 m_10 inst_913(.i1(i5[11]),
              .i2(m1200),
              .o1(m771));
 m_12 inst_914(.i1(m1195),
              .i2(m1196),
              .i3(m770),
              .o1(m772));
 m_12 inst_915(.i1(i4[12]),
              .i2(m1198),
              .i3(m772),
              .o1(m773));
 m_5 inst_916(.i1(m773),
             .o1(o17[12]));
 m_17 inst_917(.i1(i4[12]),
              .i2(m770),
              .i3(i4[13]),
              .i4(m775),
              .o1(m774));
 m_5 inst_918(.i1(i5[13]),
             .o1(m775));
 m_12 inst_919(.i1(m775),
              .i2(m1200),
              .i3(m776),
              .o1(o21[13]));
 m_10 inst_920(.i1(i5[12]),
              .i2(m1200),
              .o1(m776));
 m_12 inst_921(.i1(m1195),
              .i2(m1196),
              .i3(m775),
              .o1(m777));
 m_12 inst_922(.i1(i4[13]),
              .i2(m1198),
              .i3(m777),
              .o1(m778));
 m_5 inst_923(.i1(m778),
             .o1(o17[13]));
 m_13 inst_924(.i1(m780),
              .i2(m793),
              .i3(m798),
              .o1(m779));
 m_8 inst_925(.i1(m781),
             .i2(m790),
             .o1(m780));
 m_17 inst_926(.i1(i4[10]),
              .i2(m782),
              .i3(i4[11]),
              .i4(m786),
              .o1(m781));
 m_5 inst_927(.i1(i5[10]),
             .o1(m782));
 m_12 inst_928(.i1(m782),
              .i2(m1200),
              .i3(m783),
              .o1(o21[10]));
 m_10 inst_929(.i1(i5[9]),
              .i2(m1200),
              .o1(m783));
 m_12 inst_930(.i1(m1195),
              .i2(m1196),
              .i3(m782),
              .o1(m784));
 m_12 inst_931(.i1(i4[10]),
              .i2(m1198),
              .i3(m784),
              .o1(m785));
 m_5 inst_932(.i1(m785),
             .o1(o17[10]));
 m_5 inst_933(.i1(i5[11]),
             .o1(m786));
 m_12 inst_934(.i1(m786),
              .i2(m1200),
              .i3(m787),
              .o1(o21[11]));
 m_10 inst_935(.i1(i5[10]),
              .i2(m1200),
              .o1(m787));
 m_12 inst_936(.i1(m1195),
              .i2(m1196),
              .i3(m786),
              .o1(m788));
 m_12 inst_937(.i1(i4[11]),
              .i2(m1198),
              .i3(m788),
              .o1(m789));
 m_5 inst_938(.i1(m789),
             .o1(o17[11]));
 m_17 inst_939(.i1(m791),
              .i2(i5[10]),
              .i3(m752),
              .i4(i5[11]),
              .o1(m790));
 m_5 inst_940(.i1(i4[10]),
             .o1(m791));
 m_12 inst_941(.i1(m791),
              .i2(m185),
              .i3(m792),
              .o1(o20[11]));
 m_12 inst_942(.i1(m182),
              .i2(m183),
              .i3(i4[11]),
              .o1(m792));
 m_10 inst_943(.i1(i4[9]),
              .i2(m794),
              .o1(m793));
 m_5 inst_944(.i1(i5[9]),
             .o1(m794));
 m_12 inst_945(.i1(m794),
              .i2(m1200),
              .i3(m795),
              .o1(o21[9]));
 m_10 inst_946(.i1(i5[8]),
              .i2(m1200),
              .o1(m795));
 m_12 inst_947(.i1(m1195),
              .i2(m1196),
              .i3(m794),
              .o1(m796));
 m_12 inst_948(.i1(i4[9]),
              .i2(m1198),
              .i3(m796),
              .o1(m797));
 m_5 inst_949(.i1(m797),
             .o1(o17[9]));
 m_14 inst_950(.i1(i4[8]),
              .i2(m799),
              .i3(m803),
              .o1(m798));
 m_5 inst_951(.i1(i5[8]),
             .o1(m799));
 m_12 inst_952(.i1(m799),
              .i2(m1200),
              .i3(m800),
              .o1(o21[8]));
 m_10 inst_953(.i1(i5[7]),
              .i2(m1200),
              .o1(m800));
 m_12 inst_954(.i1(m1195),
              .i2(m1196),
              .i3(m799),
              .o1(m801));
 m_12 inst_955(.i1(i4[8]),
              .i2(m1198),
              .i3(m801),
              .o1(m802));
 m_5 inst_956(.i1(m802),
             .o1(o17[8]));
 m_17 inst_957(.i1(i4[8]),
              .i2(m799),
              .i3(i4[9]),
              .i4(m794),
              .o1(m803));
 m_12 inst_958(.i1(m804),
              .i2(m819),
              .i3(m748),
              .o1(m827));
 m_12 inst_959(.i1(m805),
              .i2(m810),
              .i3(m818),
              .o1(m804));
 m_16 inst_960(.i1(i4[6]),
              .i2(m806),
              .o1(m805));
 m_5 inst_961(.i1(i5[6]),
             .o1(m806));
 m_12 inst_962(.i1(m806),
              .i2(m1200),
              .i3(m807),
              .o1(o21[6]));
 m_10 inst_963(.i1(i5[5]),
              .i2(m1200),
              .o1(m807));
 m_12 inst_964(.i1(m1195),
              .i2(m1196),
              .i3(m806),
              .o1(m808));
 m_12 inst_965(.i1(i4[6]),
              .i2(m1198),
              .i3(m808),
              .o1(m809));
 m_5 inst_966(.i1(m809),
             .o1(o17[6]));
 m_14 inst_967(.i1(i4[5]),
              .i2(m811),
              .i3(m810),
              .o1(m884));
 m_5 inst_968(.i1(i5[5]),
             .o1(m811));
 m_12 inst_969(.i1(m811),
              .i2(m1200),
              .i3(m812),
              .o1(o21[5]));
 m_10 inst_970(.i1(i5[4]),
              .i2(m1200),
              .o1(m812));
 m_12 inst_971(.i1(m1195),
              .i2(m1196),
              .i3(m811),
              .o1(m813));
 m_12 inst_972(.i1(i4[5]),
              .i2(m1198),
              .i3(m813),
              .o1(m814));
 m_5 inst_973(.i1(m814),
             .o1(o17[5]));
 m_8 inst_974(.i1(m815),
             .i2(i5[7]),
             .o1(m810));
 m_5 inst_975(.i1(i4[7]),
             .o1(m815));
 m_12 inst_976(.i1(m815),
              .i2(m185),
              .i3(m817),
              .o1(o20[8]));
 m_12 inst_977(.i1(m815),
              .i2(m1200),
              .i3(m816),
              .o1(o20[7]));
 m_10 inst_978(.i1(i4[6]),
              .i2(m1200),
              .o1(m816));
 m_12 inst_979(.i1(m182),
              .i2(m183),
              .i3(i4[8]),
              .o1(m817));
 m_10 inst_980(.i1(m815),
              .i2(i5[7]),
              .o1(m818));
 m_14 inst_981(.i1(m820),
              .i2(m824),
              .i3(m883),
              .o1(m819));
 m_19 inst_982(.i1(m887),
              .i2(i5[4]),
              .i3(m821),
              .i4(i5[5]),
              .o1(m820));
 m_5 inst_983(.i1(i4[5]),
             .o1(m821));
 m_12 inst_984(.i1(m821),
              .i2(m185),
              .i3(m823),
              .o1(o20[6]));
 m_12 inst_985(.i1(m821),
              .i2(m1200),
              .i3(m822),
              .o1(o20[5]));
 m_10 inst_986(.i1(i4[4]),
              .i2(m1200),
              .o1(m822));
 m_12 inst_987(.i1(m182),
              .i2(m183),
              .i3(i4[6]),
              .o1(m823));
 m_12 inst_988(.i1(m887),
              .i2(i5[4]),
              .i3(m825),
              .o1(m824));
 m_12 inst_989(.i1(i4[3]),
              .i2(m857),
              .i3(m826),
              .o1(m825));
 m_13 inst_990(.i1(m827),
              .i2(m828),
              .i3(m832),
              .o1(m833));
 m_12 inst_991(.i1(m829),
              .i2(i5[15]),
              .i3(m756),
              .o1(m828));
 m_5 inst_992(.i1(i4[15]),
             .o1(m829));
 m_12 inst_993(.i1(m829),
              .i2(m185),
              .i3(m831),
              .o1(o20[16]));
 m_12 inst_994(.i1(m829),
              .i2(m1200),
              .i3(m830),
              .o1(o20[15]));
 m_10 inst_995(.i1(i4[14]),
              .i2(m1200),
              .o1(m830));
 m_12 inst_996(.i1(m182),
              .i2(m183),
              .i3(i4[16]),
              .o1(m831));
 m_14 inst_997(.i1(m889),
              .i2(m833),
              .i3(m834),
              .o1(m270));
 m_12 inst_998(.i1(m890),
              .i2(m906),
              .i3(m835),
              .o1(m834));
 m_12 inst_999(.i1(m836),
              .i2(i5[19]),
              .i3(m891),
              .o1(m835));
 m_5 inst_1000(.i1(i4[19]),
              .o1(m836));
 m_8 inst_1001(.i1(m838),
              .i2(m876),
              .o1(m837));
 m_13 inst_1002(.i1(m839),
               .i2(m855),
               .i3(m868),
               .o1(m838));
 m_5 inst_1003(.i1(m839),
              .o1(m269));
 m_8 inst_1004(.i1(m840),
              .i2(m849),
              .o1(m839));
 m_17 inst_1005(.i1(i4[20]),
               .i2(m841),
               .i3(i4[21]),
               .i4(m845),
               .o1(m840));
 m_5 inst_1006(.i1(i5[20]),
              .o1(m841));
 m_12 inst_1007(.i1(m841),
               .i2(m1200),
               .i3(m842),
               .o1(o21[20]));
 m_10 inst_1008(.i1(i5[19]),
               .i2(m1200),
               .o1(m842));
 m_12 inst_1009(.i1(m1195),
               .i2(m1196),
               .i3(m841),
               .o1(m843));
 m_12 inst_1010(.i1(i4[20]),
               .i2(m1198),
               .i3(m843),
               .o1(m844));
 m_5 inst_1011(.i1(m844),
              .o1(o17[20]));
 m_5 inst_1012(.i1(i5[21]),
              .o1(m845));
 m_12 inst_1013(.i1(m845),
               .i2(m1200),
               .i3(m846),
               .o1(o21[21]));
 m_10 inst_1014(.i1(i5[20]),
               .i2(m1200),
               .o1(m846));
 m_12 inst_1015(.i1(m1195),
               .i2(m1196),
               .i3(m845),
               .o1(m847));
 m_12 inst_1016(.i1(i4[21]),
               .i2(m1198),
               .i3(m847),
               .o1(m848));
 m_5 inst_1017(.i1(m848),
              .o1(o17[21]));
 m_17 inst_1018(.i1(m850),
               .i2(i5[20]),
               .i3(m853),
               .i4(i5[21]),
               .o1(m849));
 m_5 inst_1019(.i1(i4[20]),
              .o1(m850));
 m_12 inst_1020(.i1(m850),
               .i2(m185),
               .i3(m852),
               .o1(o20[21]));
 m_12 inst_1021(.i1(m850),
               .i2(m1200),
               .i3(m851),
               .o1(o20[20]));
 m_10 inst_1022(.i1(i4[19]),
               .i2(m1200),
               .o1(m851));
 m_12 inst_1023(.i1(m182),
               .i2(m183),
               .i3(i4[21]),
               .o1(m852));
 m_5 inst_1024(.i1(i4[21]),
              .o1(m853));
 m_12 inst_1025(.i1(m853),
               .i2(m185),
               .i3(m854),
               .o1(o20[22]));
 m_12 inst_1026(.i1(m182),
               .i2(m183),
               .i3(i4[22]),
               .o1(m854));
 m_8 inst_1027(.i1(m856),
              .i2(m867),
              .o1(m855));
 m_19 inst_1028(.i1(i4[3]),
               .i2(m857),
               .i3(m856),
               .i4(m861),
               .o1(m864));
 m_5 inst_1029(.i1(i5[3]),
              .o1(m857));
 m_12 inst_1030(.i1(m857),
               .i2(m1200),
               .i3(m858),
               .o1(o21[3]));
 m_10 inst_1031(.i1(i5[2]),
               .i2(m1200),
               .o1(m858));
 m_12 inst_1032(.i1(m1195),
               .i2(m1196),
               .i3(m857),
               .o1(m859));
 m_12 inst_1033(.i1(i4[3]),
               .i2(m1198),
               .i3(m859),
               .o1(m860));
 m_5 inst_1034(.i1(m860),
              .o1(o17[3]));
 m_19 inst_1035(.i1(m865),
               .i2(i5[1]),
               .i3(m862),
               .i4(i5[2]),
               .o1(m861));
 m_5 inst_1036(.i1(i4[2]),
              .o1(m862));
 m_12 inst_1037(.i1(m862),
               .i2(m185),
               .i3(m863),
               .o1(o20[3]));
 m_12 inst_1038(.i1(m182),
               .i2(m183),
               .i3(i4[3]),
               .o1(m863));
 m_12 inst_1039(.i1(m862),
               .i2(i5[2]),
               .i3(m864),
               .o1(m826));
 m_17 inst_1040(.i1(m879),
               .i2(i5[0]),
               .i3(m865),
               .i4(i5[1]),
               .o1(m856));
 m_5 inst_1041(.i1(i4[1]),
              .o1(m865));
 m_12 inst_1042(.i1(m865),
               .i2(m185),
               .i3(m866),
               .o1(o20[2]));
 m_12 inst_1043(.i1(m182),
               .i2(m183),
               .i3(i4[2]),
               .o1(m866));
 m_20 inst_1044(.i1(i4[2]),
               .i2(i5[2]),
               .o1(m867));
 m_8 inst_1045(.i1(m869),
              .i2(m870),
              .o1(m868));
 m_10 inst_1046(.i1(m739),
               .i2(m288),
               .o1(m869));
 m_12 inst_1047(.i1(i4[1]),
               .i2(m871),
               .i3(m875),
               .o1(m870));
 m_5 inst_1048(.i1(i5[1]),
              .o1(m871));
 m_12 inst_1049(.i1(m871),
               .i2(m1200),
               .i3(m872),
               .o1(o21[1]));
 m_10 inst_1050(.i1(i5[0]),
               .i2(m1200),
               .o1(m872));
 m_12 inst_1051(.i1(m1195),
               .i2(m1196),
               .i3(m871),
               .o1(m873));
 m_12 inst_1052(.i1(i4[1]),
               .i2(m1198),
               .i3(m873),
               .o1(m874));
 m_5 inst_1053(.i1(m874),
              .o1(o17[1]));
 m_6 inst_1054(.i1(i4[3]),
              .i2(i5[3]),
              .o1(m875));
 m_10 inst_1055(.i1(m877),
               .i2(m878),
               .o1(m876));
 m_14 inst_1056(.i1(m879),
               .i2(i5[0]),
               .i3(m311),
               .o1(m878));
 m_5 inst_1057(.i1(i4[0]),
              .o1(m879));
 m_8 inst_1058(.i1(m879),
              .i2(m1200),
              .o1(o20[0]));
 m_12 inst_1059(.i1(m879),
               .i2(m185),
               .i3(m880),
               .o1(o20[1]));
 m_12 inst_1060(.i1(m182),
               .i2(m183),
               .i3(i4[1]),
               .o1(m880));
 m_8 inst_1061(.i1(m882),
              .i2(m888),
              .o1(m881));
 m_16 inst_1062(.i1(m883),
               .i2(m886),
               .o1(m882));
 m_13 inst_1063(.i1(m818),
               .i2(m884),
               .i3(m885),
               .o1(m883));
 m_6 inst_1064(.i1(i4[6]),
              .i2(i5[6]),
              .o1(m885));
 m_12 inst_1065(.i1(m887),
               .i2(i5[4]),
               .i3(m820),
               .o1(m886));
 m_5 inst_1066(.i1(i4[4]),
              .o1(m887));
 m_13 inst_1067(.i1(m889),
               .i2(m907),
               .i3(m908),
               .o1(m888));
 m_8 inst_1068(.i1(m890),
              .i2(m903),
              .o1(m889));
 m_16 inst_1069(.i1(m891),
               .i2(m900),
               .o1(m890));
 m_17 inst_1070(.i1(i4[18]),
               .i2(m892),
               .i3(i4[19]),
               .i4(m896),
               .o1(m891));
 m_5 inst_1071(.i1(i5[18]),
              .o1(m892));
 m_12 inst_1072(.i1(m892),
               .i2(m1200),
               .i3(m893),
               .o1(o21[18]));
 m_10 inst_1073(.i1(i5[17]),
               .i2(m1200),
               .o1(m893));
 m_12 inst_1074(.i1(m1195),
               .i2(m1196),
               .i3(m892),
               .o1(m894));
 m_12 inst_1075(.i1(i4[18]),
               .i2(m1198),
               .i3(m894),
               .o1(m895));
 m_5 inst_1076(.i1(m895),
              .o1(o17[18]));
 m_5 inst_1077(.i1(i5[19]),
              .o1(m896));
 m_12 inst_1078(.i1(m896),
               .i2(m1200),
               .i3(m897),
               .o1(o21[19]));
 m_10 inst_1079(.i1(i5[18]),
               .i2(m1200),
               .o1(m897));
 m_12 inst_1080(.i1(m1195),
               .i2(m1196),
               .i3(m896),
               .o1(m898));
 m_12 inst_1081(.i1(i4[19]),
               .i2(m1198),
               .i3(m898),
               .o1(m899));
 m_5 inst_1082(.i1(m899),
              .o1(o17[19]));
 m_12 inst_1083(.i1(m901),
               .i2(i5[17]),
               .i3(m902),
               .o1(m900));
 m_5 inst_1084(.i1(i4[17]),
              .o1(m901));
 m_19 inst_1085(.i1(i4[18]),
               .i2(m892),
               .i3(i4[19]),
               .i4(m896),
               .o1(m902));
 m_12 inst_1086(.i1(m904),
               .i2(i5[16]),
               .i3(m906),
               .o1(m903));
 m_5 inst_1087(.i1(i4[16]),
              .o1(m904));
 m_12 inst_1088(.i1(m904),
               .i2(m185),
               .i3(m905),
               .o1(o20[17]));
 m_12 inst_1089(.i1(m182),
               .i2(m183),
               .i3(i4[17]),
               .o1(m905));
 m_19 inst_1090(.i1(m904),
               .i2(i5[16]),
               .i3(m901),
               .i4(i5[17]),
               .o1(m906));
 m_6 inst_1091(.i1(i4[22]),
              .i2(i5[22]),
              .o1(m907));
 m_8 inst_1092(.i1(m185),
              .i2(m909),
              .o1(m908));
 m_6 inst_1093(.i1(i3[0]),
              .i2(m909),
              .o1(o13));
 m_20 inst_1094(.i1(i4[31]),
               .i2(i5[31]),
               .o1(m909));
 m_13 inst_1095(.i1(m910),
               .i2(m1023),
               .i3(m1108),
               .o1(o16));
 m_18 inst_1096(.i1(i4[31]),
               .i2(m910),
               .i3(m911),
               .o1(m914));
 m_10 inst_1097(.i1(o14[1]),
               .i2(m912),
               .o1(m911));
 m_15 inst_1098(.i1(o14[1]),
               .i2(m912),
               .o1(m913));
 m_8 inst_1099(.i1(i3[3]),
              .i2(i3[2]),
              .o1(m912));
 m_14 inst_1100(.i1(m915),
               .i2(m917),
               .i3(m914),
               .o1(m922));
 m_12 inst_1101(.i1(o14[1]),
               .i2(m916),
               .i3(i3[3]),
               .o1(m915));
 m_13 inst_1102(.i1(m928),
               .i2(m919),
               .i3(m920),
               .o1(m916));
 m_14 inst_1103(.i1(m918),
               .i2(m913),
               .i3(m921),
               .o1(m917));
 m_13 inst_1104(.i1(m919),
               .i2(m920),
               .i3(m1117),
               .o1(m918));
 m_16 inst_1105(.i1(m925),
               .i2(m926),
               .o1(m919));
 m_12 inst_1106(.i1(m925),
               .i2(m926),
               .i3(m920),
               .o1(o14[0]));
 m_5 inst_1107(.i1(i4[31]),
              .o1(m921));
 m_14 inst_1108(.i1(m922),
               .i2(m1178),
               .i3(m923),
               .o1(o3[0]));
 m_12 inst_1109(.i1(m922),
               .i2(m1178),
               .i3(m1321),
               .o1(m923));
 m_18 inst_1110(.i1(m924),
               .i2(m933),
               .i3(m969),
               .o1(m910));
 m_8 inst_1111(.i1(m925),
              .i2(m926),
              .o1(m924));
 m_18 inst_1112(.i1(m924),
               .i2(m933),
               .i3(o14[1]),
               .o1(m927));
 m_14 inst_1113(.i1(m928),
               .i2(m927),
               .i3(m932),
               .o1(m1020));
 m_15 inst_1114(.i1(i3[1]),
               .i2(m928),
               .o1(m929));
 m_12 inst_1115(.i1(m1208),
               .i2(m930),
               .i3(m931),
               .o1(m928));
 m_10 inst_1116(.i1(i4[29]),
               .i2(i4[28]),
               .o1(m930));
 m_5 inst_1117(.i1(i4[30]),
              .o1(m931));
 m_5 inst_1118(.i1(i3[3]),
              .o1(m932));
 m_13 inst_1119(.i1(m934),
               .i2(m939),
               .i3(m946),
               .o1(m933));
 m_12 inst_1120(.i1(m935),
               .i2(m971),
               .i3(m938),
               .o1(m934));
 m_2 inst_1121(.i1(m1007),
              .i2(m936),
              .i3(m945),
              .o1(m935));
 m_2 inst_1122(.i1(m1015),
              .i2(m937),
              .i3(m943),
              .o1(m936));
 m_8 inst_1123(.i1(m243),
              .i2(m977),
              .o1(m937));
 m_5 inst_1124(.i1(m938),
              .o1(m989));
 m_12 inst_1125(.i1(m940),
               .i2(m944),
               .i3(m945),
               .o1(m939));
 m_2 inst_1126(.i1(m941),
              .i2(m942),
              .i3(m943),
              .o1(m940));
 m_2 inst_1127(.i1(m1153),
              .i2(m1132),
              .i3(m257),
              .o1(m941));
 m_2 inst_1128(.i1(m1155),
              .i2(m1138),
              .i3(m257),
              .o1(m942));
 m_13 inst_1129(.i1(m936),
               .i2(m1000),
               .i3(m975),
               .o1(m944));
 m_8 inst_1130(.i1(m947),
              .i2(m963),
              .o1(m946));
 m_14 inst_1131(.i1(m948),
               .i2(m949),
               .i3(m243),
               .o1(m947));
 m_12 inst_1132(.i1(m240),
               .i2(m929),
               .i3(m1319),
               .o1(m948));
 m_12 inst_1133(.i1(m950),
               .i2(m954),
               .i3(m958),
               .o1(m949));
 m_10 inst_1134(.i1(m951),
               .i2(m857),
               .o1(m950));
 m_5 inst_1135(.i1(i5[0]),
              .o1(m951));
 m_8 inst_1136(.i1(m951),
              .i2(m1200),
              .o1(o21[0]));
 m_12 inst_1137(.i1(m1195),
               .i2(m1196),
               .i3(m951),
               .o1(m952));
 m_12 inst_1138(.i1(i4[0]),
               .i2(m1198),
               .i3(m952),
               .o1(m953));
 m_5 inst_1139(.i1(m953),
              .o1(o17[0]));
 m_13 inst_1140(.i1(m955),
               .i2(m956),
               .i3(m957),
               .o1(m954));
 m_8 inst_1141(.i1(i5[5]),
              .i2(i5[6]),
              .o1(m955));
 m_8 inst_1142(.i1(i5[4]),
              .i2(i5[7]),
              .o1(m956));
 m_8 inst_1143(.i1(i5[1]),
              .i2(i5[2]),
              .o1(m957));
 m_8 inst_1144(.i1(i3[1]),
              .i2(m1198),
              .o1(m958));
 m_16 inst_1145(.i1(m947),
               .i2(m963),
               .o1(m959));
 m_18 inst_1146(.i1(m960),
               .i2(m961),
               .i3(m959),
               .o1(m920));
 m_14 inst_1147(.i1(m962),
               .i2(m1145),
               .i3(m988),
               .o1(m961));
 m_14 inst_1148(.i1(m964),
               .i2(m966),
               .i3(m968),
               .o1(m963));
 m_18 inst_1149(.i1(m1012),
               .i2(m986),
               .i3(m965),
               .o1(m964));
 m_18 inst_1150(.i1(m1001),
               .i2(m980),
               .i3(m967),
               .o1(m966));
 m_12 inst_1151(.i1(m243),
               .i2(m1005),
               .i3(m977),
               .o1(m967));
 m_5 inst_1152(.i1(m943),
              .o1(m968));
 m_2 inst_1153(.i1(m970),
              .i2(m990),
              .i3(m925),
              .o1(m969));
 m_2 inst_1154(.i1(m926),
              .i2(m970),
              .i3(m925),
              .o1(o14[1]));
 m_2 inst_1155(.i1(m971),
              .i2(m978),
              .i3(m989),
              .o1(m970));
 m_2 inst_1156(.i1(m972),
              .i2(m975),
              .i3(m945),
              .o1(m971));
 m_2 inst_1157(.i1(m973),
              .i2(m974),
              .i3(m943),
              .o1(m972));
 m_2 inst_1158(.i1(m1009),
              .i2(m997),
              .i3(m243),
              .o1(m973));
 m_10 inst_1159(.i1(m968),
               .i2(m973),
               .o1(m1071));
 m_12 inst_1160(.i1(m243),
               .i2(m258),
               .i3(m254),
               .o1(m974));
 m_2 inst_1161(.i1(m1035),
              .i2(m976),
              .i3(m943),
              .o1(m975));
 m_2 inst_1162(.i1(m977),
              .i2(m1005),
              .i3(m243),
              .o1(m976));
 m_2 inst_1163(.i1(m979),
              .i2(m981),
              .i3(m988),
              .o1(m978));
 m_2 inst_1164(.i1(m1074),
              .i2(m980),
              .i3(m943),
              .o1(m979));
 m_2 inst_1165(.i1(m249),
              .i2(m1002),
              .i3(m257),
              .o1(m980));
 m_2 inst_1166(.i1(m982),
              .i2(m986),
              .i3(m943),
              .o1(m981));
 m_2 inst_1167(.i1(m994),
              .i2(m983),
              .i3(m243),
              .o1(m982));
 m_15 inst_1168(.i1(m984),
               .i2(m985),
               .o1(m983));
 m_13 inst_1169(.i1(m1454),
               .i2(i2[1]),
               .i3(m314),
               .o1(m984));
 m_12 inst_1170(.i1(m240),
               .i2(m929),
               .i3(i2[0]),
               .o1(m985));
 m_10 inst_1171(.i1(m968),
               .i2(m982),
               .o1(m1073));
 m_12 inst_1172(.i1(m243),
               .i2(m1016),
               .i3(m987),
               .o1(m986));
 m_12 inst_1173(.i1(m255),
               .i2(m256),
               .i3(m252),
               .o1(m987));
 m_5 inst_1174(.i1(m945),
              .o1(m988));
 m_2 inst_1175(.i1(m991),
              .i2(m1006),
              .i3(m989),
              .o1(m990));
 m_2 inst_1176(.i1(m935),
              .i2(m991),
              .i3(m989),
              .o1(m926));
 m_2 inst_1177(.i1(m992),
              .i2(m1000),
              .i3(m945),
              .o1(m991));
 m_2 inst_1178(.i1(m993),
              .i2(m999),
              .i3(m943),
              .o1(m992));
 m_2 inst_1179(.i1(m994),
              .i2(m997),
              .i3(m257),
              .o1(m993));
 m_17 inst_1180(.i1(i4[22]),
               .i2(m314),
               .i3(m240),
               .i4(m995),
               .o1(m994));
 m_12 inst_1181(.i1(i3[1]),
               .i2(m262),
               .i3(m996),
               .o1(m995));
 m_10 inst_1182(.i1(i4[22]),
               .i2(m929),
               .o1(m996));
 m_12 inst_1183(.i1(i4[21]),
               .i2(m314),
               .i3(m998),
               .o1(m997));
 m_12 inst_1184(.i1(i3[1]),
               .i2(m314),
               .i3(m1124),
               .o1(m998));
 m_10 inst_1185(.i1(m968),
               .i2(m993),
               .o1(m1028));
 m_2 inst_1186(.i1(m1029),
              .i2(m1001),
              .i3(m943),
              .o1(m1000));
 m_2 inst_1187(.i1(m1002),
              .i2(m1005),
              .i3(m257),
              .o1(m1001));
 m_17 inst_1188(.i1(i4[10]),
               .i2(m314),
               .i3(m240),
               .i4(m1003),
               .o1(m1002));
 m_12 inst_1189(.i1(i3[1]),
               .i2(m782),
               .i3(m1004),
               .o1(m1003));
 m_10 inst_1190(.i1(i4[10]),
               .i2(m929),
               .o1(m1004));
 m_2 inst_1191(.i1(m1007),
              .i2(m1013),
              .i3(m988),
              .o1(m1006));
 m_2 inst_1192(.i1(m1008),
              .i2(m1012),
              .i3(m943),
              .o1(m1007));
 m_2 inst_1193(.i1(m1009),
              .i2(m1075),
              .i3(m257),
              .o1(m1008));
 m_17 inst_1194(.i1(i4[20]),
               .i2(m314),
               .i3(m240),
               .i4(m1010),
               .o1(m1009));
 m_12 inst_1195(.i1(i3[1]),
               .i2(m841),
               .i3(m1011),
               .o1(m1010));
 m_10 inst_1196(.i1(i4[20]),
               .i2(m929),
               .o1(m1011));
 m_2 inst_1197(.i1(m1014),
              .i2(m1015),
              .i3(m943),
              .o1(m1013));
 m_10 inst_1198(.i1(m968),
               .i2(m1014),
               .o1(m1296));
 m_8 inst_1199(.i1(m257),
              .i2(m983),
              .o1(m1014));
 m_2 inst_1200(.i1(m1036),
              .i2(m1016),
              .i3(m257),
              .o1(m1015));
 m_17 inst_1201(.i1(i4[15]),
               .i2(m314),
               .i3(m240),
               .i4(m1017),
               .o1(m1016));
 m_12 inst_1202(.i1(i3[1]),
               .i2(m761),
               .i3(m1018),
               .o1(m1017));
 m_10 inst_1203(.i1(i4[15]),
               .i2(m929),
               .o1(m1018));
 m_12 inst_1204(.i1(m910),
               .i2(m911),
               .i3(i4[31]),
               .o1(m1019));
 m_12 inst_1205(.i1(m1020),
               .i2(m1019),
               .i3(m1021),
               .o1(m1022));
 m_13 inst_1206(.i1(m921),
               .i2(m918),
               .i3(m913),
               .o1(m1021));
 m_8 inst_1207(.i1(m1024),
              .i2(m1089),
              .o1(m1023));
 m_2 inst_1208(.i1(m1025),
              .i2(m1032),
              .i3(m925),
              .o1(m1024));
 m_12 inst_1209(.i1(m989),
               .i2(m1026),
               .i3(m1031),
               .o1(m1025));
 m_12 inst_1210(.i1(m988),
               .i2(m1027),
               .i3(m1030),
               .o1(m1026));
 m_2 inst_1211(.i1(m1028),
              .i2(m1027),
              .i3(m945),
              .o1(m1096));
 m_10 inst_1212(.i1(m968),
               .i2(m1029),
               .o1(m1027));
 m_2 inst_1213(.i1(m1079),
              .i2(m1044),
              .i3(m257),
              .o1(m1029));
 m_10 inst_1214(.i1(m988),
               .i2(m1119),
               .o1(m1030));
 m_10 inst_1215(.i1(m989),
               .i2(m1146),
               .o1(m1031));
 m_2 inst_1216(.i1(m1033),
              .i2(m1065),
              .i3(m989),
              .o1(m1032));
 m_12 inst_1217(.i1(m988),
               .i2(m1034),
               .i3(m1052),
               .o1(m1033));
 m_10 inst_1218(.i1(m968),
               .i2(m1035),
               .o1(m1034));
 m_2 inst_1219(.i1(m1036),
              .i2(m1044),
              .i3(m243),
              .o1(m1035));
 m_17 inst_1220(.i1(i4[16]),
               .i2(m314),
               .i3(m240),
               .i4(m1037),
               .o1(m1036));
 m_8 inst_1221(.i1(m240),
              .i2(m1037),
              .o1(m1038));
 m_12 inst_1222(.i1(i3[1]),
               .i2(m1039),
               .i3(m1043),
               .o1(m1037));
 m_5 inst_1223(.i1(i5[16]),
              .o1(m1039));
 m_12 inst_1224(.i1(m1039),
               .i2(m1200),
               .i3(m1040),
               .o1(o21[16]));
 m_10 inst_1225(.i1(i5[15]),
               .i2(m1200),
               .o1(m1040));
 m_12 inst_1226(.i1(m1195),
               .i2(m1196),
               .i3(m1039),
               .o1(m1041));
 m_12 inst_1227(.i1(i4[16]),
               .i2(m1198),
               .i3(m1041),
               .o1(m1042));
 m_5 inst_1228(.i1(m1042),
              .o1(o17[16]));
 m_10 inst_1229(.i1(i4[16]),
               .i2(m929),
               .o1(m1043));
 m_17 inst_1230(.i1(i4[17]),
               .i2(m314),
               .i3(m240),
               .i4(m1045),
               .o1(m1044));
 m_8 inst_1231(.i1(m240),
              .i2(m1045),
              .o1(m1046));
 m_12 inst_1232(.i1(i3[1]),
               .i2(m1047),
               .i3(m1051),
               .o1(m1045));
 m_5 inst_1233(.i1(i5[17]),
              .o1(m1047));
 m_12 inst_1234(.i1(m1047),
               .i2(m1200),
               .i3(m1048),
               .o1(o21[17]));
 m_10 inst_1235(.i1(i5[16]),
               .i2(m1200),
               .o1(m1048));
 m_12 inst_1236(.i1(m1195),
               .i2(m1196),
               .i3(m1047),
               .o1(m1049));
 m_12 inst_1237(.i1(i4[17]),
               .i2(m1198),
               .i3(m1049),
               .o1(m1050));
 m_5 inst_1238(.i1(m1050),
              .o1(o17[17]));
 m_10 inst_1239(.i1(i4[17]),
               .i2(m929),
               .o1(m1051));
 m_10 inst_1240(.i1(m988),
               .i2(m1053),
               .o1(m1052));
 m_2 inst_1241(.i1(m1053),
              .i2(m1054),
              .i3(m945),
              .o1(m1116));
 m_2 inst_1242(.i1(m1055),
              .i2(m1056),
              .i3(m943),
              .o1(m1054));
 m_2 inst_1243(.i1(m1161),
              .i2(m1136),
              .i3(m243),
              .o1(m1055));
 m_2 inst_1244(.i1(m1057),
              .i2(m1140),
              .i3(m243),
              .o1(m1056));
 m_14 inst_1245(.i1(m1058),
               .i2(m1198),
               .i3(m1060),
               .o1(m1057));
 m_5 inst_1246(.i1(i4[8]),
              .o1(m1058));
 m_12 inst_1247(.i1(m1058),
               .i2(m185),
               .i3(m1059),
               .o1(o20[9]));
 m_12 inst_1248(.i1(m182),
               .i2(m183),
               .i3(i4[9]),
               .o1(m1059));
 m_8 inst_1249(.i1(m240),
              .i2(m1061),
              .o1(m1060));
 m_12 inst_1250(.i1(i3[1]),
               .i2(m799),
               .i3(m1062),
               .o1(m1061));
 m_10 inst_1251(.i1(i4[8]),
               .i2(m929),
               .o1(m1062));
 m_17 inst_1252(.i1(i4[8]),
               .i2(m314),
               .i3(m240),
               .i4(m1061),
               .o1(m977));
 m_2 inst_1253(.i1(m1063),
              .i2(m1064),
              .i3(m943),
              .o1(m1053));
 m_2 inst_1254(.i1(m1151),
              .i2(m1123),
              .i3(m243),
              .o1(m1063));
 m_2 inst_1255(.i1(m244),
              .i2(m1126),
              .i3(m243),
              .o1(m1064));
 m_2 inst_1256(.i1(m1066),
              .i2(m1065),
              .i3(m938),
              .o1(m1094));
 m_2 inst_1257(.i1(m1067),
              .i2(m1066),
              .i3(m938),
              .o1(m1070));
 m_12 inst_1258(.i1(m938),
               .i2(m1067),
               .i3(m1068),
               .o1(m1069));
 m_12 inst_1259(.i1(m945),
               .i2(m1071),
               .i3(m938),
               .o1(m1068));
 m_2 inst_1260(.i1(m1099),
              .i2(m1069),
              .i3(m1293),
              .o1(o14[7]));
 m_2 inst_1261(.i1(m1103),
              .i2(m1070),
              .i3(m1293),
              .o1(o14[5]));
 m_2 inst_1262(.i1(m1071),
              .i2(m1034),
              .i3(m945),
              .o1(m1066));
 m_12 inst_1263(.i1(m945),
               .i2(m1071),
               .i3(m989),
               .o1(m1101));
 m_12 inst_1264(.i1(m988),
               .i2(m1072),
               .i3(m1083),
               .o1(m1065));
 m_2 inst_1265(.i1(m1073),
              .i2(m1072),
              .i3(m945),
              .o1(m1067));
 m_12 inst_1266(.i1(m945),
               .i2(m1073),
               .i3(m938),
               .o1(m1102));
 m_10 inst_1267(.i1(m968),
               .i2(m1074),
               .o1(m1072));
 m_2 inst_1268(.i1(m1075),
              .i2(m1079),
              .i3(m257),
              .o1(m1074));
 m_17 inst_1269(.i1(i4[19]),
               .i2(m314),
               .i3(m240),
               .i4(m1076),
               .o1(m1075));
 m_8 inst_1270(.i1(m240),
              .i2(m1076),
              .o1(m1077));
 m_12 inst_1271(.i1(i3[1]),
               .i2(m896),
               .i3(m1078),
               .o1(m1076));
 m_10 inst_1272(.i1(i4[19]),
               .i2(m929),
               .o1(m1078));
 m_17 inst_1273(.i1(i4[18]),
               .i2(m314),
               .i3(m240),
               .i4(m1080),
               .o1(m1079));
 m_8 inst_1274(.i1(m240),
              .i2(m1080),
              .o1(m1081));
 m_12 inst_1275(.i1(i3[1]),
               .i2(m892),
               .i3(m1082),
               .o1(m1080));
 m_10 inst_1276(.i1(i4[18]),
               .i2(m929),
               .o1(m1082));
 m_10 inst_1277(.i1(m988),
               .i2(m1084),
               .o1(m1083));
 m_2 inst_1278(.i1(m1085),
              .i2(m1087),
              .i3(m943),
              .o1(m1084));
 m_2 inst_1279(.i1(m1121),
              .i2(m1086),
              .i3(m243),
              .o1(m1085));
 m_10 inst_1280(.i1(m984),
               .i2(m985),
               .o1(m1086));
 m_2 inst_1281(.i1(m1162),
              .i2(m252),
              .i3(m257),
              .o1(m1087));
 m_6 inst_1282(.i1(i4[31]),
              .i2(m1024),
              .o1(m1088));
 m_16 inst_1283(.i1(m1090),
               .i2(m1092),
               .o1(m1089));
 m_2 inst_1284(.i1(m1110),
              .i2(m1025),
              .i3(m925),
              .o1(m1090));
 m_6 inst_1285(.i1(i4[31]),
              .i2(m1090),
              .o1(m1091));
 m_2 inst_1286(.i1(m1032),
              .i2(m1093),
              .i3(m925),
              .o1(m1092));
 m_2 inst_1287(.i1(m1093),
              .i2(m1094),
              .i3(m925),
              .o1(o14[2]));
 m_2 inst_1288(.i1(m1094),
              .i2(m1104),
              .i3(m925),
              .o1(o14[3]));
 m_2 inst_1289(.i1(m1026),
              .i2(m1095),
              .i3(m989),
              .o1(m1093));
 m_2 inst_1290(.i1(m1096),
              .i2(m1095),
              .i3(m938),
              .o1(m1104));
 m_2 inst_1291(.i1(m1097),
              .i2(m1096),
              .i3(m938),
              .o1(m1103));
 m_12 inst_1292(.i1(m938),
               .i2(m1097),
               .i3(m1098),
               .o1(m1099));
 m_12 inst_1293(.i1(m945),
               .i2(m1028),
               .i3(m938),
               .o1(m1098));
 m_2 inst_1294(.i1(m1100),
              .i2(m1099),
              .i3(m1293),
              .o1(o14[8]));
 m_10 inst_1295(.i1(m1101),
               .i2(m1102),
               .o1(m1100));
 m_2 inst_1296(.i1(m1103),
              .i2(m1069),
              .i3(m925),
              .o1(o14[6]));
 m_2 inst_1297(.i1(m1070),
              .i2(m1104),
              .i3(m1293),
              .o1(o14[4]));
 m_12 inst_1298(.i1(m988),
               .i2(m1105),
               .i3(m1106),
               .o1(m1095));
 m_2 inst_1299(.i1(m1296),
              .i2(m1105),
              .i3(m945),
              .o1(m1097));
 m_10 inst_1300(.i1(m968),
               .i2(m1008),
               .o1(m1105));
 m_10 inst_1301(.i1(m988),
               .i2(m1157),
               .o1(m1106));
 m_6 inst_1302(.i1(i4[31]),
              .i2(m1092),
              .o1(m1107));
 m_8 inst_1303(.i1(o14[1]),
              .i2(m1109),
              .o1(m1108));
 m_12 inst_1304(.i1(m925),
               .i2(m1110),
               .i3(m1113),
               .o1(m1109));
 m_12 inst_1305(.i1(m989),
               .i2(m1033),
               .i3(m1111),
               .o1(m1110));
 m_10 inst_1306(.i1(m989),
               .i2(m1112),
               .o1(m1111));
 m_2 inst_1307(.i1(m940),
              .i2(m1084),
              .i3(m988),
              .o1(m1112));
 m_10 inst_1308(.i1(m925),
               .i2(m1114),
               .o1(m1113));
 m_2 inst_1309(.i1(m1115),
              .i2(m1114),
              .i3(m925),
              .o1(m1117));
 m_2 inst_1310(.i1(m1116),
              .i2(m1112),
              .i3(m989),
              .o1(m1115));
 m_14 inst_1311(.i1(m1149),
               .i2(m1116),
               .i3(m989),
               .o1(m960));
 m_2 inst_1312(.i1(m1118),
              .i2(m1146),
              .i3(m989),
              .o1(m1114));
 m_2 inst_1313(.i1(m1119),
              .i2(m1130),
              .i3(m945),
              .o1(m1118));
 m_2 inst_1314(.i1(m1120),
              .i2(m1125),
              .i3(m943),
              .o1(m1119));
 m_2 inst_1315(.i1(m1121),
              .i2(m1123),
              .i3(m257),
              .o1(m1120));
 m_14 inst_1316(.i1(m267),
               .i2(m1198),
               .i3(m1122),
               .o1(m1121));
 m_8 inst_1317(.i1(m240),
              .i2(m995),
              .o1(m1122));
 m_19 inst_1318(.i1(m853),
               .i2(m1198),
               .i3(m276),
               .i4(m1124),
               .o1(m1123));
 m_19 inst_1319(.i1(m1454),
               .i2(i5[21]),
               .i3(m929),
               .i4(i4[21]),
               .o1(m1124));
 m_2 inst_1320(.i1(m252),
              .i2(m1126),
              .i3(m257),
              .o1(m1125));
 m_14 inst_1321(.i1(m766),
               .i2(m1198),
               .i3(m1127),
               .o1(m1126));
 m_8 inst_1322(.i1(m240),
              .i2(m1128),
              .o1(m1127));
 m_12 inst_1323(.i1(i3[1]),
               .i2(m775),
               .i3(m1129),
               .o1(m1128));
 m_10 inst_1324(.i1(i4[13]),
               .i2(m929),
               .o1(m1129));
 m_2 inst_1325(.i1(m1131),
              .i2(m1137),
              .i3(m943),
              .o1(m1130));
 m_2 inst_1326(.i1(m1132),
              .i2(m1136),
              .i3(m257),
              .o1(m1131));
 m_14 inst_1327(.i1(m1133),
               .i2(m1198),
               .i3(m1081),
               .o1(m1132));
 m_5 inst_1328(.i1(i4[18]),
              .o1(m1133));
 m_12 inst_1329(.i1(m1133),
               .i2(m185),
               .i3(m1135),
               .o1(o20[19]));
 m_12 inst_1330(.i1(m1133),
               .i2(m1200),
               .i3(m1134),
               .o1(o20[18]));
 m_10 inst_1331(.i1(i4[17]),
               .i2(m1200),
               .o1(m1134));
 m_12 inst_1332(.i1(m182),
               .i2(m183),
               .i3(i4[19]),
               .o1(m1135));
 m_14 inst_1333(.i1(m901),
               .i2(m1198),
               .i3(m1046),
               .o1(m1136));
 m_2 inst_1334(.i1(m1138),
              .i2(m1140),
              .i3(m257),
              .o1(m1137));
 m_14 inst_1335(.i1(m791),
               .i2(m1198),
               .i3(m1139),
               .o1(m1138));
 m_8 inst_1336(.i1(m240),
              .i2(m1003),
              .o1(m1139));
 m_19 inst_1337(.i1(m1141),
               .i2(m1198),
               .i3(m276),
               .i4(m1143),
               .o1(m1140));
 m_5 inst_1338(.i1(i4[9]),
              .o1(m1141));
 m_12 inst_1339(.i1(m1141),
               .i2(m185),
               .i3(m1142),
               .o1(o20[10]));
 m_12 inst_1340(.i1(m182),
               .i2(m183),
               .i3(i4[10]),
               .o1(m1142));
 m_19 inst_1341(.i1(m1454),
               .i2(i5[9]),
               .i3(m929),
               .i4(i4[9]),
               .o1(m1143));
 m_12 inst_1342(.i1(i3[1]),
               .i2(m314),
               .i3(m1143),
               .o1(m1144));
 m_12 inst_1343(.i1(i4[9]),
               .i2(m314),
               .i3(m1144),
               .o1(m1005));
 m_8 inst_1344(.i1(m1130),
              .i2(m940),
              .o1(m1145));
 m_2 inst_1345(.i1(m1147),
              .i2(m1157),
              .i3(m988),
              .o1(m1146));
 m_2 inst_1346(.i1(m1147),
              .i2(m1148),
              .i3(m945),
              .o1(m1149));
 m_8 inst_1347(.i1(m1148),
              .i2(m1054),
              .o1(m962));
 m_2 inst_1348(.i1(m1150),
              .i2(m1154),
              .i3(m943),
              .o1(m1147));
 m_2 inst_1349(.i1(m1151),
              .i2(m1153),
              .i3(m257),
              .o1(m1150));
 m_14 inst_1350(.i1(m850),
               .i2(m1198),
               .i3(m1152),
               .o1(m1151));
 m_8 inst_1351(.i1(m240),
              .i2(m1010),
              .o1(m1152));
 m_14 inst_1352(.i1(m836),
               .i2(m1198),
               .i3(m1077),
               .o1(m1153));
 m_2 inst_1353(.i1(m244),
              .i2(m1155),
              .i3(m257),
              .o1(m1154));
 m_14 inst_1354(.i1(m752),
               .i2(m1198),
               .i3(m1156),
               .o1(m1155));
 m_2 inst_1355(.i1(m1158),
              .i2(m1159),
              .i3(m943),
              .o1(m1157));
 m_12 inst_1356(.i1(m255),
               .i2(m256),
               .i3(m1086),
               .o1(m1158));
 m_2 inst_1357(.i1(m1159),
              .i2(m1160),
              .i3(m943),
              .o1(m1148));
 m_10 inst_1358(.i1(m257),
               .i2(m1057),
               .o1(m1160));
 m_2 inst_1359(.i1(m1161),
              .i2(m1162),
              .i3(m257),
              .o1(m1159));
 m_14 inst_1360(.i1(m904),
               .i2(m1198),
               .i3(m1038),
               .o1(m1161));
 m_14 inst_1361(.i1(m829),
               .i2(m1198),
               .i3(m1163),
               .o1(m1162));
 m_8 inst_1362(.i1(m240),
              .i2(m1017),
              .o1(m1163));
 m_6 inst_1363(.i1(i4[31]),
              .i2(m1109),
              .o1(m1164));
 m_5 inst_1364(.i1(m1164),
              .o1(m1165));
 m_13 inst_1365(.i1(m1022),
               .i2(m1166),
               .i3(m1165),
               .o1(m1167));
 m_5 inst_1366(.i1(m1166),
              .o1(m1178));
 m_6 inst_1367(.i1(i4[31]),
              .i2(m1117),
              .o1(m1166));
 m_14 inst_1368(.i1(m1167),
               .i2(m1091),
               .i3(m1173),
               .o1(o3[2]));
 m_18 inst_1369(.i1(m1167),
               .i2(m1091),
               .i3(m1088),
               .o1(m1168));
 m_10 inst_1370(.i1(m1168),
               .i2(m1169),
               .o1(m1170));
 m_5 inst_1371(.i1(m1107),
              .o1(m1169));
 m_14 inst_1372(.i1(m1170),
               .i2(m1247),
               .i3(m1171),
               .o1(o3[5]));
 m_12 inst_1373(.i1(m1170),
               .i2(m1247),
               .i3(m1321),
               .o1(m1171));
 m_13 inst_1374(.i1(m1168),
               .i2(m1169),
               .i3(m1172),
               .o1(m1241));
 m_5 inst_1375(.i1(m1247),
              .o1(m1172));
 m_12 inst_1376(.i1(m1167),
               .i2(m1091),
               .i3(m1321),
               .o1(m1173));
 m_12 inst_1377(.i1(m1174),
               .i2(m1165),
               .i3(m1175),
               .o1(m1177));
 m_8 inst_1378(.i1(m922),
              .i2(m1178),
              .o1(m1174));
 m_8 inst_1379(.i1(m1179),
              .i2(m1176),
              .o1(m1175));
 m_5 inst_1380(.i1(m1321),
              .o1(m1176));
 m_5 inst_1381(.i1(m1177),
              .o1(o3[1]));
 m_18 inst_1382(.i1(m922),
               .i2(m1178),
               .i3(m1164),
               .o1(m1179));
 m_10 inst_1383(.i1(m1179),
               .i2(m1180),
               .o1(m1181));
 m_5 inst_1384(.i1(m1091),
              .o1(m1180));
 m_14 inst_1385(.i1(m1181),
               .i2(m1088),
               .i3(m1182),
               .o1(o3[3]));
 m_12 inst_1386(.i1(m1181),
               .i2(m1088),
               .i3(m1321),
               .o1(m1182));
 m_13 inst_1387(.i1(m1179),
               .i2(m1180),
               .i3(m1183),
               .o1(m1184));
 m_5 inst_1388(.i1(m1088),
              .o1(m1183));
 m_14 inst_1389(.i1(m1184),
               .i2(m1107),
               .i3(m1185),
               .o1(o3[4]));
 m_12 inst_1390(.i1(m1184),
               .i2(m1107),
               .i3(m1321),
               .o1(m1185));
 m_5 inst_1391(.i1(m620),
              .o1(o19));
 m_12 inst_1392(.i1(m1194),
               .i2(m1200),
               .i3(m1201),
               .o1(o21[7]));
 m_12 inst_1393(.i1(m1186),
               .i2(m1200),
               .i3(m1189),
               .o1(o21[4]));
 m_5 inst_1394(.i1(i5[4]),
              .o1(m1186));
 m_12 inst_1395(.i1(m1195),
               .i2(m1196),
               .i3(m1186),
               .o1(m1187));
 m_12 inst_1396(.i1(i4[4]),
               .i2(m1198),
               .i3(m1187),
               .o1(m1188));
 m_5 inst_1397(.i1(m1188),
              .o1(o17[4]));
 m_10 inst_1398(.i1(i5[3]),
               .i2(m1200),
               .o1(m1189));
 m_12 inst_1399(.i1(m1190),
               .i2(m1200),
               .i3(m1193),
               .o1(o21[2]));
 m_5 inst_1400(.i1(i5[2]),
              .o1(m1190));
 m_12 inst_1401(.i1(m1195),
               .i2(m1196),
               .i3(m1190),
               .o1(m1191));
 m_12 inst_1402(.i1(i4[2]),
               .i2(m1198),
               .i3(m1191),
               .o1(m1192));
 m_5 inst_1403(.i1(m1192),
              .o1(o17[2]));
 m_10 inst_1404(.i1(i5[1]),
               .i2(m1200),
               .o1(m1193));
 m_5 inst_1405(.i1(i5[7]),
              .o1(m1194));
 m_12 inst_1406(.i1(m1195),
               .i2(m1196),
               .i3(m1194),
               .o1(m1197));
 m_12 inst_1407(.i1(i4[7]),
               .i2(m1198),
               .i3(m1197),
               .o1(m1199));
 m_5 inst_1408(.i1(m1199),
              .o1(o17[7]));
 m_10 inst_1409(.i1(i5[6]),
               .i2(m1200),
               .o1(m1201));
 m_14 inst_1410(.i1(m1202),
               .i2(m1204),
               .i3(o15),
               .o1(o2));
 m_16 inst_1411(.i1(i4[31]),
               .i2(m1203),
               .o1(m1202));
 m_10 inst_1412(.i1(i5[31]),
               .i2(m1203),
               .o1(m1204));
 m_12 inst_1413(.i1(m1203),
               .i2(m1205),
               .i3(m1204),
               .o1(o6[33]));
 m_6 inst_1414(.i1(i4[31]),
              .i2(i3[0]),
              .o1(m1205));
 m_14 inst_1415(.i1(m1206),
               .i2(m1262),
               .i3(m1318),
               .o1(o7));
 m_19 inst_1416(.i1(i4[30]),
               .i2(m1207),
               .i3(m1237),
               .i4(m1261),
               .o1(m1206));
 m_13 inst_1417(.i1(m1208),
               .i2(m1209),
               .i3(m1212),
               .o1(m1207));
 m_12 inst_1418(.i1(i4[27]),
               .i2(m1210),
               .i3(m1211),
               .o1(m1209));
 m_10 inst_1419(.i1(i4[27]),
               .i2(m1210),
               .o1(m1208));
 m_14 inst_1420(.i1(m659),
               .i2(m705),
               .i3(i1[1]),
               .o1(m1211));
 m_5 inst_1421(.i1(m1213),
              .o1(m1212));
 m_12 inst_1422(.i1(m1214),
               .i2(m1218),
               .i3(m1219),
               .o1(m1213));
 m_8 inst_1423(.i1(i4[26]),
              .i2(m1215),
              .o1(m1214));
 m_15 inst_1424(.i1(i4[26]),
               .i2(m1215),
               .o1(m1210));
 m_8 inst_1425(.i1(m742),
              .i2(m703),
              .o1(m1215));
 m_12 inst_1426(.i1(m1210),
               .i2(m1214),
               .i3(i3[1]),
               .o1(m1216));
 m_12 inst_1427(.i1(i3[1]),
               .i2(m1217),
               .i3(m1216),
               .o1(m943));
 m_17 inst_1428(.i1(m295),
               .i2(m745),
               .i3(m237),
               .i4(m236),
               .o1(m1217));
 m_12 inst_1429(.i1(i4[26]),
               .i2(i4[23]),
               .i3(m1261),
               .o1(m1218));
 m_13 inst_1430(.i1(i4[30]),
               .i2(m1219),
               .i3(m1220),
               .o1(m1224));
 m_8 inst_1431(.i1(i4[23]),
              .i2(m1221),
              .o1(m1220));
 m_10 inst_1432(.i1(m267),
               .i2(i1[1]),
               .o1(m1221));
 m_12 inst_1433(.i1(i4[31]),
               .i2(m1221),
               .i3(m1222),
               .o1(m1223));
 m_14 inst_1434(.i1(i4[22]),
               .i2(i4[31]),
               .i3(m1302),
               .o1(m1222));
 m_5 inst_1435(.i1(m1223),
              .o1(m547));
 m_8 inst_1436(.i1(m1208),
              .i2(m1224),
              .o1(m1225));
 m_13 inst_1437(.i1(m1225),
               .i2(m1226),
               .i3(m1230),
               .o1(m1320));
 m_8 inst_1438(.i1(m1227),
              .i2(m1228),
              .o1(m1226));
 m_13 inst_1439(.i1(m850),
               .i2(m853),
               .i3(i4[31]),
               .o1(m1227));
 m_13 inst_1440(.i1(m1133),
               .i2(m836),
               .i3(m1229),
               .o1(m1228));
 m_8 inst_1441(.i1(i4[16]),
              .i2(i4[17]),
              .o1(m1229));
 m_15 inst_1442(.i1(m752),
               .i2(m1231),
               .o1(m1230));
 m_8 inst_1443(.i1(m1232),
              .i2(m1236),
              .o1(m1231));
 m_13 inst_1444(.i1(m1233),
               .i2(m829),
               .i3(m1235),
               .o1(m1232));
 m_19 inst_1445(.i1(m1233),
               .i2(m1198),
               .i3(m276),
               .i4(m1234),
               .o1(m252));
 m_19 inst_1446(.i1(m1454),
               .i2(i5[14]),
               .i3(m929),
               .i4(i4[14]),
               .o1(m1234));
 m_5 inst_1447(.i1(i4[14]),
              .o1(m1233));
 m_8 inst_1448(.i1(i4[12]),
              .i2(i4[13]),
              .o1(m1235));
 m_13 inst_1449(.i1(m1058),
               .i2(m1141),
               .i3(m791),
               .o1(m1236));
 m_8 inst_1450(.i1(i4[29]),
              .i2(i4[28]),
              .o1(m1219));
 m_6 inst_1451(.i1(m1238),
              .i2(m1239),
              .o1(m1237));
 m_12 inst_1452(.i1(m1319),
               .i2(m1320),
               .i3(m1239),
               .o1(m1240));
 m_8 inst_1453(.i1(m1253),
              .i2(m1240),
              .o1(o3[7]));
 m_12 inst_1454(.i1(m1241),
               .i2(m1243),
               .i3(m1244),
               .o1(m1239));
 m_14 inst_1455(.i1(m1241),
               .i2(m1243),
               .i3(m1242),
               .o1(o3[6]));
 m_12 inst_1456(.i1(m1241),
               .i2(m1243),
               .i3(m1321),
               .o1(m1242));
 m_6 inst_1457(.i1(i4[31]),
              .i2(o14[3]),
              .o1(m1243));
 m_5 inst_1458(.i1(m1244),
              .o1(m1245));
 m_13 inst_1459(.i1(m1246),
               .i2(m1248),
               .i3(m1245),
               .o1(m1249));
 m_18 inst_1460(.i1(m1184),
               .i2(m1107),
               .i3(m1247),
               .o1(m1246));
 m_6 inst_1461(.i1(i4[31]),
              .i2(o14[2]),
              .o1(m1247));
 m_5 inst_1462(.i1(m1243),
              .o1(m1248));
 m_14 inst_1463(.i1(m1238),
               .i2(m1249),
               .i3(m1252),
               .o1(o3[8]));
 m_18 inst_1464(.i1(m1238),
               .i2(m1249),
               .i3(m1258),
               .o1(m1250));
 m_13 inst_1465(.i1(m1250),
               .i2(m1251),
               .i3(m1273),
               .o1(m1265));
 m_5 inst_1466(.i1(m1271),
              .o1(m1251));
 m_12 inst_1467(.i1(m1238),
               .i2(m1249),
               .i3(m1321),
               .o1(m1252));
 m_18 inst_1468(.i1(m1241),
               .i2(m1243),
               .i3(m1244),
               .o1(m1253));
 m_10 inst_1469(.i1(m1254),
               .i2(m1253),
               .o1(m1255));
 m_5 inst_1470(.i1(m1254),
              .o1(m1238));
 m_6 inst_1471(.i1(m921),
              .i2(o14[5]),
              .o1(m1254));
 m_14 inst_1472(.i1(m1255),
               .i2(m1258),
               .i3(m1256),
               .o1(o3[9]));
 m_12 inst_1473(.i1(m1255),
               .i2(m1258),
               .i3(m1321),
               .o1(m1256));
 m_13 inst_1474(.i1(m1254),
               .i2(m1253),
               .i3(m1257),
               .o1(m1259));
 m_5 inst_1475(.i1(m1258),
              .o1(m1257));
 m_6 inst_1476(.i1(i4[31]),
              .i2(o14[6]),
              .o1(m1258));
 m_14 inst_1477(.i1(m1259),
               .i2(m1271),
               .i3(m1260),
               .o1(o3[10]));
 m_12 inst_1478(.i1(m1259),
               .i2(m1271),
               .i3(m1321),
               .o1(m1260));
 m_6 inst_1479(.i1(i4[31]),
              .i2(o14[4]),
              .o1(m1244));
 m_8 inst_1480(.i1(i1[1]),
              .i2(i1[0]),
              .o1(m1261));
 m_13 inst_1481(.i1(m1263),
               .i2(m1298),
               .i3(m1310),
               .o1(m1262));
 m_13 inst_1482(.i1(m1264),
               .i2(m1280),
               .i3(m1292),
               .o1(m1263));
 m_18 inst_1483(.i1(m1265),
               .i2(m1267),
               .i3(m1268),
               .o1(m1264));
 m_14 inst_1484(.i1(m1265),
               .i2(m1267),
               .i3(m1266),
               .o1(o3[12]));
 m_12 inst_1485(.i1(m1265),
               .i2(m1267),
               .i3(m1321),
               .o1(m1266));
 m_14 inst_1486(.i1(m1278),
               .i2(m1268),
               .i3(m1279),
               .o1(o3[13]));
 m_5 inst_1487(.i1(m1269),
              .o1(m1268));
 m_13 inst_1488(.i1(m1270),
               .i2(m1277),
               .i3(m1269),
               .o1(m1311));
 m_18 inst_1489(.i1(m1259),
               .i2(m1271),
               .i3(m1272),
               .o1(m1270));
 m_6 inst_1490(.i1(i4[31]),
              .i2(o14[7]),
              .o1(m1271));
 m_5 inst_1491(.i1(m1273),
              .o1(m1272));
 m_8 inst_1492(.i1(m1274),
              .i2(m1273),
              .o1(m1275));
 m_8 inst_1493(.i1(m1259),
              .i2(m1271),
              .o1(m1274));
 m_8 inst_1494(.i1(m1275),
              .i2(m1276),
              .o1(o3[11]));
 m_12 inst_1495(.i1(m1319),
               .i2(m1320),
               .i3(m1265),
               .o1(m1276));
 m_6 inst_1496(.i1(m921),
              .i2(o14[8]),
              .o1(m1273));
 m_5 inst_1497(.i1(m1267),
              .o1(m1277));
 m_6 inst_1498(.i1(i4[31]),
              .i2(m1290),
              .o1(m1269));
 m_12 inst_1499(.i1(m1278),
               .i2(m1268),
               .i3(m1321),
               .o1(m1279));
 m_10 inst_1500(.i1(m1270),
               .i2(m1277),
               .o1(m1278));
 m_5 inst_1501(.i1(m1280),
              .o1(m1316));
 m_6 inst_1502(.i1(i4[31]),
              .i2(m1281),
              .o1(m1280));
 m_14 inst_1503(.i1(m925),
               .i2(m1282),
               .i3(m1291),
               .o1(m1281));
 m_8 inst_1504(.i1(m938),
              .i2(m1283),
              .o1(m1282));
 m_12 inst_1505(.i1(m938),
               .i2(m1283),
               .i3(m1293),
               .o1(m1284));
 m_12 inst_1506(.i1(m1293),
               .i2(m1285),
               .i3(m1284),
               .o1(m1290));
 m_15 inst_1507(.i1(m1286),
               .i2(m1287),
               .o1(m1285));
 m_12 inst_1508(.i1(m945),
               .i2(m1028),
               .i3(m989),
               .o1(m1286));
 m_12 inst_1509(.i1(m945),
               .i2(m1296),
               .i3(m938),
               .o1(m1287));
 m_12 inst_1510(.i1(m925),
               .i2(m1285),
               .i3(m1288),
               .o1(m1289));
 m_10 inst_1511(.i1(m925),
               .i2(m1100),
               .o1(m1288));
 m_5 inst_1512(.i1(m1289),
              .o1(o14[9]));
 m_6 inst_1513(.i1(m921),
              .i2(m1289),
              .o1(m1267));
 m_5 inst_1514(.i1(m1290),
              .o1(o14[10]));
 m_16 inst_1515(.i1(m945),
               .i2(m1073),
               .o1(m1283));
 m_8 inst_1516(.i1(m925),
              .i2(m1294),
              .o1(m1291));
 m_5 inst_1517(.i1(m1281),
              .o1(o14[11]));
 m_12 inst_1518(.i1(m1293),
               .i2(m1294),
               .i3(m921),
               .o1(m1292));
 m_5 inst_1519(.i1(m1293),
              .o1(m925));
 m_10 inst_1520(.i1(m989),
               .i2(m1295),
               .o1(m1294));
 m_8 inst_1521(.i1(m945),
              .i2(m1296),
              .o1(m1295));
 m_8 inst_1522(.i1(m1293),
              .i2(m1294),
              .o1(o14[12]));
 m_12 inst_1523(.i1(o14[12]),
               .i2(m1263),
               .i3(i4[31]),
               .o1(m1297));
 m_8 inst_1524(.i1(m1297),
              .i2(m1176),
              .o1(o3[18]));
 m_8 inst_1525(.i1(m1297),
              .i2(m1176),
              .o1(o3[17]));
 m_8 inst_1526(.i1(m1297),
              .i2(m1176),
              .o1(o3[16]));
 m_12 inst_1527(.i1(m1319),
               .i2(m1320),
               .i3(m1297),
               .o1(o3[19]));
 m_8 inst_1528(.i1(i1[1]),
              .i2(m1299),
              .o1(m1298));
 m_5 inst_1529(.i1(i1[0]),
              .o1(m1299));
 m_18 inst_1530(.i1(i4[15]),
               .i2(i1[1]),
               .i3(m1299),
               .o1(m1300));
 m_18 inst_1531(.i1(m1301),
               .i2(m1303),
               .i3(m1300),
               .o1(m1309));
 m_8 inst_1532(.i1(m1302),
              .i2(i4[31]),
              .o1(m1301));
 m_5 inst_1533(.i1(i1[1]),
              .o1(m1302));
 m_8 inst_1534(.i1(i4[7]),
              .i2(m1304),
              .o1(m1303));
 m_12 inst_1535(.i1(i4[7]),
               .i2(m1304),
               .i3(m1305),
               .o1(m232));
 m_5 inst_1536(.i1(m614),
              .o1(m1305));
 m_17 inst_1537(.i1(m815),
               .i2(m1304),
               .i3(m1306),
               .i4(m829),
               .o1(m1308));
 m_10 inst_1538(.i1(m1302),
               .i2(i1[0]),
               .o1(m1306));
 m_12 inst_1539(.i1(i4[15]),
               .i2(m1306),
               .i3(m1307),
               .o1(m614));
 m_10 inst_1540(.i1(i1[1]),
               .i2(m921),
               .o1(m1307));
 m_16 inst_1541(.i1(i1[1]),
               .i2(i1[0]),
               .o1(m1304));
 m_12 inst_1542(.i1(m1311),
               .i2(m1316),
               .i3(m1317),
               .o1(m1310));
 m_14 inst_1543(.i1(m1311),
               .i2(m1316),
               .i3(m1315),
               .o1(o3[14]));
 m_8 inst_1544(.i1(m1311),
              .i2(m1316),
              .o1(m1312));
 m_14 inst_1545(.i1(m1312),
               .i2(m1313),
               .i3(m1314),
               .o1(o3[15]));
 m_12 inst_1546(.i1(m1312),
               .i2(m1313),
               .i3(m1321),
               .o1(m1314));
 m_6 inst_1547(.i1(m921),
              .i2(o14[12]),
              .o1(m1313));
 m_12 inst_1548(.i1(m1311),
               .i2(m1316),
               .i3(m1321),
               .o1(m1315));
 m_5 inst_1549(.i1(o14[12]),
              .o1(m1317));
 m_12 inst_1550(.i1(m1319),
               .i2(m1320),
               .i3(m1322),
               .o1(m1318));
 m_16 inst_1551(.i1(m1319),
               .i2(m1320),
               .o1(m1321));
 m_15 inst_1552(.i1(i3[1]),
               .i2(i3[0]),
               .o1(m1322));
 m_8 inst_1553(.i1(i3[1]),
              .i2(m1323),
              .o1(o8));
 m_14 inst_1554(.i1(m1323),
               .i2(m1324),
               .i3(m1325),
               .o1(o6[0]));
 m_14 inst_1555(.i1(i18[1]),
               .i2(i18[26]),
               .i3(i18[0]),
               .o1(m1324));
 m_14 inst_1556(.i1(i18[2]),
               .i2(m1326),
               .i3(m1394),
               .o1(m1325));
 m_12 inst_1557(.i1(i18[25]),
               .i2(m1326),
               .i3(o13),
               .o1(m1393));
 m_12 inst_1558(.i1(i18[24]),
               .i2(m1326),
               .i3(m1357),
               .o1(m1358));
 m_12 inst_1559(.i1(i18[15]),
               .i2(m1326),
               .i3(m1327),
               .o1(m1328));
 m_5 inst_1560(.i1(m1425),
              .o1(m1327));
 m_12 inst_1561(.i1(o13),
               .i2(m1329),
               .i3(m1328),
               .o1(o6[14]));
 m_2 inst_1562(.i1(i18[15]),
              .i2(i18[14]),
              .i3(i18[26]),
              .o1(m1329));
 m_12 inst_1563(.i1(i18[14]),
               .i2(m1326),
               .i3(m1330),
               .o1(m1331));
 m_5 inst_1564(.i1(m1426),
              .o1(m1330));
 m_12 inst_1565(.i1(o13),
               .i2(m1332),
               .i3(m1331),
               .o1(o6[13]));
 m_2 inst_1566(.i1(i18[14]),
              .i2(i18[13]),
              .i3(i18[26]),
              .o1(m1332));
 m_12 inst_1567(.i1(i18[13]),
               .i2(m1326),
               .i3(m1333),
               .o1(m1334));
 m_5 inst_1568(.i1(m1427),
              .o1(m1333));
 m_12 inst_1569(.i1(o13),
               .i2(m1335),
               .i3(m1334),
               .o1(o6[12]));
 m_2 inst_1570(.i1(i18[13]),
              .i2(i18[12]),
              .i3(i18[26]),
              .o1(m1335));
 m_12 inst_1571(.i1(i18[12]),
               .i2(m1326),
               .i3(m1336),
               .o1(m1337));
 m_5 inst_1572(.i1(m1428),
              .o1(m1336));
 m_12 inst_1573(.i1(o13),
               .i2(m1338),
               .i3(m1337),
               .o1(o6[11]));
 m_2 inst_1574(.i1(i18[12]),
              .i2(i18[11]),
              .i3(i18[26]),
              .o1(m1338));
 m_12 inst_1575(.i1(i18[11]),
               .i2(m1326),
               .i3(m1339),
               .o1(m1340));
 m_5 inst_1576(.i1(m1429),
              .o1(m1339));
 m_12 inst_1577(.i1(o13),
               .i2(m1341),
               .i3(m1340),
               .o1(o6[10]));
 m_2 inst_1578(.i1(i18[11]),
              .i2(i18[10]),
              .i3(i18[26]),
              .o1(m1341));
 m_12 inst_1579(.i1(i18[10]),
               .i2(m1326),
               .i3(m1342),
               .o1(m1343));
 m_5 inst_1580(.i1(m1430),
              .o1(m1342));
 m_12 inst_1581(.i1(o13),
               .i2(m1344),
               .i3(m1343),
               .o1(o6[9]));
 m_2 inst_1582(.i1(i18[10]),
              .i2(i18[9]),
              .i3(i18[26]),
              .o1(m1344));
 m_12 inst_1583(.i1(i18[9]),
               .i2(m1326),
               .i3(m1345),
               .o1(m1346));
 m_5 inst_1584(.i1(m1431),
              .o1(m1345));
 m_12 inst_1585(.i1(o13),
               .i2(m1347),
               .i3(m1346),
               .o1(o6[8]));
 m_2 inst_1586(.i1(i18[9]),
              .i2(i18[8]),
              .i3(i18[26]),
              .o1(m1347));
 m_12 inst_1587(.i1(i18[8]),
               .i2(m1326),
               .i3(m1348),
               .o1(m1349));
 m_5 inst_1588(.i1(m1432),
              .o1(m1348));
 m_12 inst_1589(.i1(o13),
               .i2(m1350),
               .i3(m1349),
               .o1(o6[7]));
 m_2 inst_1590(.i1(i18[8]),
              .i2(i18[7]),
              .i3(i18[26]),
              .o1(m1350));
 m_12 inst_1591(.i1(i18[7]),
               .i2(m1326),
               .i3(m1351),
               .o1(m1352));
 m_5 inst_1592(.i1(m1433),
              .o1(m1351));
 m_12 inst_1593(.i1(o13),
               .i2(m1353),
               .i3(m1352),
               .o1(o6[6]));
 m_2 inst_1594(.i1(i18[7]),
              .i2(i18[6]),
              .i3(i18[26]),
              .o1(m1353));
 m_12 inst_1595(.i1(i18[6]),
               .i2(m1326),
               .i3(m1354),
               .o1(m1355));
 m_5 inst_1596(.i1(m1434),
              .o1(m1354));
 m_12 inst_1597(.i1(o13),
               .i2(m1356),
               .i3(m1355),
               .o1(o6[5]));
 m_2 inst_1598(.i1(i18[6]),
              .i2(i18[5]),
              .i3(i18[26]),
              .o1(m1356));
 m_5 inst_1599(.i1(m1435),
              .o1(m1357));
 m_12 inst_1600(.i1(o13),
               .i2(m1359),
               .i3(m1358),
               .o1(o6[23]));
 m_2 inst_1601(.i1(i18[24]),
              .i2(i18[23]),
              .i3(i18[26]),
              .o1(m1359));
 m_12 inst_1602(.i1(i18[23]),
               .i2(m1326),
               .i3(m1369),
               .o1(m1370));
 m_12 inst_1603(.i1(i18[5]),
               .i2(m1326),
               .i3(m1360),
               .o1(m1361));
 m_5 inst_1604(.i1(m1436),
              .o1(m1360));
 m_12 inst_1605(.i1(o13),
               .i2(m1362),
               .i3(m1361),
               .o1(o6[4]));
 m_2 inst_1606(.i1(i18[5]),
              .i2(i18[4]),
              .i3(i18[26]),
              .o1(m1362));
 m_12 inst_1607(.i1(i18[4]),
               .i2(m1326),
               .i3(m1363),
               .o1(m1364));
 m_5 inst_1608(.i1(m1437),
              .o1(m1363));
 m_12 inst_1609(.i1(o13),
               .i2(m1365),
               .i3(m1364),
               .o1(o6[3]));
 m_2 inst_1610(.i1(i18[4]),
              .i2(i18[3]),
              .i3(i18[26]),
              .o1(m1365));
 m_12 inst_1611(.i1(i18[2]),
               .i2(m1326),
               .i3(m1366),
               .o1(m1367));
 m_5 inst_1612(.i1(m1438),
              .o1(m1366));
 m_12 inst_1613(.i1(o13),
               .i2(m1368),
               .i3(m1367),
               .o1(o6[1]));
 m_2 inst_1614(.i1(i18[2]),
              .i2(i18[1]),
              .i3(i18[26]),
              .o1(m1368));
 m_5 inst_1615(.i1(m1439),
              .o1(m1369));
 m_12 inst_1616(.i1(o13),
               .i2(m1371),
               .i3(m1370),
               .o1(o6[22]));
 m_2 inst_1617(.i1(i18[23]),
              .i2(i18[22]),
              .i3(i18[26]),
              .o1(m1371));
 m_12 inst_1618(.i1(i18[22]),
               .i2(m1326),
               .i3(m1372),
               .o1(m1373));
 m_5 inst_1619(.i1(m1440),
              .o1(m1372));
 m_12 inst_1620(.i1(o13),
               .i2(m1374),
               .i3(m1373),
               .o1(o6[21]));
 m_2 inst_1621(.i1(i18[22]),
              .i2(i18[21]),
              .i3(i18[26]),
              .o1(m1374));
 m_12 inst_1622(.i1(i18[21]),
               .i2(m1326),
               .i3(m1375),
               .o1(m1376));
 m_5 inst_1623(.i1(m1441),
              .o1(m1375));
 m_12 inst_1624(.i1(o13),
               .i2(m1377),
               .i3(m1376),
               .o1(o6[20]));
 m_2 inst_1625(.i1(i18[21]),
              .i2(i18[20]),
              .i3(i18[26]),
              .o1(m1377));
 m_12 inst_1626(.i1(i18[20]),
               .i2(m1326),
               .i3(m1378),
               .o1(m1379));
 m_5 inst_1627(.i1(m1442),
              .o1(m1378));
 m_12 inst_1628(.i1(o13),
               .i2(m1380),
               .i3(m1379),
               .o1(o6[19]));
 m_2 inst_1629(.i1(i18[20]),
              .i2(i18[19]),
              .i3(i18[26]),
              .o1(m1380));
 m_12 inst_1630(.i1(i18[19]),
               .i2(m1326),
               .i3(m1381),
               .o1(m1382));
 m_5 inst_1631(.i1(m1443),
              .o1(m1381));
 m_12 inst_1632(.i1(o13),
               .i2(m1383),
               .i3(m1382),
               .o1(o6[18]));
 m_2 inst_1633(.i1(i18[19]),
              .i2(i18[18]),
              .i3(i18[26]),
              .o1(m1383));
 m_12 inst_1634(.i1(i18[18]),
               .i2(m1326),
               .i3(m1384),
               .o1(m1385));
 m_5 inst_1635(.i1(m1444),
              .o1(m1384));
 m_12 inst_1636(.i1(o13),
               .i2(m1386),
               .i3(m1385),
               .o1(o6[17]));
 m_2 inst_1637(.i1(i18[18]),
              .i2(i18[17]),
              .i3(i18[26]),
              .o1(m1386));
 m_12 inst_1638(.i1(i18[17]),
               .i2(m1326),
               .i3(m1387),
               .o1(m1388));
 m_5 inst_1639(.i1(m1445),
              .o1(m1387));
 m_12 inst_1640(.i1(o13),
               .i2(m1389),
               .i3(m1388),
               .o1(o6[16]));
 m_2 inst_1641(.i1(i18[17]),
              .i2(i18[16]),
              .i3(i18[26]),
              .o1(m1389));
 m_12 inst_1642(.i1(i18[16]),
               .i2(m1326),
               .i3(m1390),
               .o1(m1391));
 m_5 inst_1643(.i1(m1446),
              .o1(m1390));
 m_12 inst_1644(.i1(o13),
               .i2(m1392),
               .i3(m1391),
               .o1(o6[15]));
 m_2 inst_1645(.i1(i18[16]),
              .i2(i18[15]),
              .i3(i18[26]),
              .o1(m1392));
 m_5 inst_1646(.i1(m1393),
              .o1(m1447));
 m_10 inst_1647(.i1(o13),
               .i2(m1395),
               .o1(m1394));
 m_8 inst_1648(.i1(i18[1]),
              .i2(i18[0]),
              .o1(m1395));
 m_5 inst_1649(.i1(o13),
              .o1(m1323));
 m_12 inst_1650(.i1(m1396),
               .i2(i18[3]),
               .i3(m1323),
               .o1(m1397));
 m_5 inst_1651(.i1(i18[26]),
              .o1(m1396));
 m_12 inst_1652(.i1(m1398),
               .i2(m1397),
               .i3(m1421),
               .o1(o6[2]));
 m_10 inst_1653(.i1(m1395),
               .i2(m1398),
               .o1(m1399));
 m_8 inst_1654(.i1(m1400),
              .i2(m1399),
              .o1(m1403));
 m_10 inst_1655(.i1(m1401),
               .i2(m1402),
               .o1(m1400));
 m_8 inst_1656(.i1(i18[3]),
              .i2(i18[4]),
              .o1(m1401));
 m_8 inst_1657(.i1(i18[5]),
              .i2(i18[6]),
              .o1(m1402));
 m_13 inst_1658(.i1(m1404),
               .i2(m1403),
               .i3(m1413),
               .o1(m1420));
 m_8 inst_1659(.i1(m1405),
              .i2(m1409),
              .o1(m1404));
 m_13 inst_1660(.i1(m1406),
               .i2(m1407),
               .i3(m1408),
               .o1(m1405));
 m_8 inst_1661(.i1(i18[20]),
              .i2(i18[21]),
              .o1(m1406));
 m_8 inst_1662(.i1(i18[19]),
              .i2(i18[22]),
              .o1(m1407));
 m_8 inst_1663(.i1(i18[15]),
              .i2(i18[18]),
              .o1(m1408));
 m_13 inst_1664(.i1(m1410),
               .i2(m1411),
               .i3(m1412),
               .o1(m1409));
 m_5 inst_1665(.i1(i18[24]),
              .o1(m1410));
 m_8 inst_1666(.i1(i18[23]),
              .i2(i18[25]),
              .o1(m1411));
 m_8 inst_1667(.i1(i18[16]),
              .i2(i18[17]),
              .o1(m1412));
 m_8 inst_1668(.i1(m1414),
              .i2(m1417),
              .o1(m1413));
 m_10 inst_1669(.i1(m1415),
               .i2(m1416),
               .o1(m1414));
 m_8 inst_1670(.i1(i18[11]),
              .i2(i18[12]),
              .o1(m1415));
 m_8 inst_1671(.i1(i18[13]),
              .i2(i18[14]),
              .o1(m1416));
 m_10 inst_1672(.i1(m1418),
               .i2(m1419),
               .o1(m1417));
 m_8 inst_1673(.i1(i18[7]),
              .i2(i18[8]),
              .o1(m1418));
 m_8 inst_1674(.i1(i18[9]),
              .i2(i18[10]),
              .o1(m1419));
 m_8 inst_1675(.i1(o13),
              .i2(m1420),
              .o1(o6[34]));
 m_8 inst_1676(.i1(i18[2]),
              .i2(i18[26]),
              .o1(m1398));
 m_12 inst_1677(.i1(i18[3]),
               .i2(m1326),
               .i3(m1422),
               .o1(m1421));
 m_5 inst_1678(.i1(m1423),
              .o1(m1422));
 m_12 inst_1679(.i1(i18[4]),
               .i2(m1424),
               .i3(o13),
               .o1(m1423));
 m_12 inst_1680(.i1(i18[26]),
               .i2(m1424),
               .i3(m1447),
               .o1(m1448));
 m_12 inst_1681(.i1(i18[25]),
               .i2(m1424),
               .i3(o13),
               .o1(m1435));
 m_12 inst_1682(.i1(i18[16]),
               .i2(m1424),
               .i3(o13),
               .o1(m1425));
 m_12 inst_1683(.i1(i18[15]),
               .i2(m1424),
               .i3(o13),
               .o1(m1426));
 m_12 inst_1684(.i1(i18[14]),
               .i2(m1424),
               .i3(o13),
               .o1(m1427));
 m_12 inst_1685(.i1(i18[13]),
               .i2(m1424),
               .i3(o13),
               .o1(m1428));
 m_12 inst_1686(.i1(i18[12]),
               .i2(m1424),
               .i3(o13),
               .o1(m1429));
 m_12 inst_1687(.i1(i18[11]),
               .i2(m1424),
               .i3(o13),
               .o1(m1430));
 m_12 inst_1688(.i1(i18[10]),
               .i2(m1424),
               .i3(o13),
               .o1(m1431));
 m_12 inst_1689(.i1(i18[9]),
               .i2(m1424),
               .i3(o13),
               .o1(m1432));
 m_12 inst_1690(.i1(i18[8]),
               .i2(m1424),
               .i3(o13),
               .o1(m1433));
 m_12 inst_1691(.i1(i18[7]),
               .i2(m1424),
               .i3(o13),
               .o1(m1434));
 m_12 inst_1692(.i1(i18[24]),
               .i2(m1424),
               .i3(o13),
               .o1(m1439));
 m_12 inst_1693(.i1(i18[6]),
               .i2(m1424),
               .i3(o13),
               .o1(m1436));
 m_12 inst_1694(.i1(i18[5]),
               .i2(m1424),
               .i3(o13),
               .o1(m1437));
 m_12 inst_1695(.i1(i18[3]),
               .i2(m1424),
               .i3(o13),
               .o1(m1438));
 m_12 inst_1696(.i1(i18[23]),
               .i2(m1424),
               .i3(o13),
               .o1(m1440));
 m_12 inst_1697(.i1(i18[22]),
               .i2(m1424),
               .i3(o13),
               .o1(m1441));
 m_12 inst_1698(.i1(i18[21]),
               .i2(m1424),
               .i3(o13),
               .o1(m1442));
 m_12 inst_1699(.i1(i18[20]),
               .i2(m1424),
               .i3(o13),
               .o1(m1443));
 m_12 inst_1700(.i1(i18[19]),
               .i2(m1424),
               .i3(o13),
               .o1(m1444));
 m_12 inst_1701(.i1(i18[18]),
               .i2(m1424),
               .i3(o13),
               .o1(m1445));
 m_12 inst_1702(.i1(i18[17]),
               .i2(m1424),
               .i3(o13),
               .o1(m1446));
 m_12 inst_1703(.i1(o13),
               .i2(m1449),
               .i3(m1448),
               .o1(o6[24]));
 m_2 inst_1704(.i1(i18[25]),
              .i2(i18[24]),
              .i3(i18[26]),
              .o1(m1449));
 m_10 inst_1705(.i1(m1454),
               .i2(m1455),
               .o1(o9[7]));
 m_10 inst_1706(.i1(m1454),
               .i2(m1450),
               .o1(o9[4]));
 m_5 inst_1707(.i1(m1450),
              .o1(o4[29]));
 m_2 inst_1708(.i1(i10[31]),
              .i2(i11[31]),
              .i3(m1203),
              .o1(m1450));
 m_10 inst_1709(.i1(m1454),
               .i2(m1451),
               .o1(o9[3]));
 m_5 inst_1710(.i1(m1451),
              .o1(o4[28]));
 m_2 inst_1711(.i1(i10[30]),
              .i2(i11[30]),
              .i3(m1203),
              .o1(m1451));
 m_10 inst_1712(.i1(m1454),
               .i2(m1452),
               .o1(o9[2]));
 m_5 inst_1713(.i1(m1452),
              .o1(o4[27]));
 m_2 inst_1714(.i1(i10[29]),
              .i2(i11[29]),
              .i3(m1203),
              .o1(m1452));
 m_10 inst_1715(.i1(m1454),
               .i2(m1453),
               .o1(o9[1]));
 m_5 inst_1716(.i1(m1453),
              .o1(o4[26]));
 m_2 inst_1717(.i1(i10[28]),
              .i2(i11[28]),
              .i3(m1203),
              .o1(m1453));
 m_5 inst_1718(.i1(i3[1]),
              .o1(m1454));
 m_5 inst_1719(.i1(m1455),
              .o1(o4[32]));
 m_2 inst_1720(.i1(i10[34]),
              .i2(i11[34]),
              .i3(m1203),
              .o1(m1455));
 m_8 inst_1721(.i1(i3[1]),
              .i2(m1460),
              .o1(o9[8]));
 m_8 inst_1722(.i1(i3[1]),
              .i2(m1456),
              .o1(o9[6]));
 m_5 inst_1723(.i1(m1456),
              .o1(o4[31]));
 m_2 inst_1724(.i1(i10[33]),
              .i2(i11[33]),
              .i3(m1203),
              .o1(m1456));
 m_8 inst_1725(.i1(i3[1]),
              .i2(m1457),
              .o1(o9[5]));
 m_5 inst_1726(.i1(m1457),
              .o1(o4[30]));
 m_2 inst_1727(.i1(i10[32]),
              .i2(i11[32]),
              .i3(m1203),
              .o1(m1457));
 m_8 inst_1728(.i1(i3[1]),
              .i2(m1458),
              .o1(o9[0]));
 m_5 inst_1729(.i1(m1458),
              .o1(o4[25]));
 m_2 inst_1730(.i1(i10[27]),
              .i2(i11[27]),
              .i3(m1203),
              .o1(m1458));
 m_6 inst_1731(.i1(m691),
              .i2(m1458),
              .o1(m1459));
 m_5 inst_1732(.i1(m1460),
              .o1(o4[33]));
 m_2 inst_1733(.i1(i10[35]),
              .i2(i11[35]),
              .i3(m1203),
              .o1(m1460));
 endmodule

 module m_20 (
    input i1,
    input i2,
    output o1
 );
 m_7 inst_1(.i1(i1),
           .i2(i2),
           .o1(o1));
 endmodule

 module m_19 (
    input i1,
    input i2,
    input i3,
    input i4,
    output o1
 );
 wire m1;
 wire m2;
 wire m3;
 m_3 inst_1(.i1(m2),
           .o1(o1));
 m_9 inst_2(.i1(m3),
           .i2(m1),
           .o1(m2));
 m_11 inst_3(.i1(i3),
            .i2(i4),
            .o1(m1));
 m_11 inst_4(.i1(i1),
            .i2(i2),
            .o1(m3));
 endmodule

 module m_18 (
    input i1,
    input i2,
    input i3,
    output o1
 );
 wire m1;
 wire m2;
 m_3 inst_1(.i1(m2),
           .o1(o1));
 m_9 inst_2(.i1(m1),
           .i2(i3),
           .o1(m2));
 m_9 inst_3(.i1(i1),
           .i2(i2),
           .o1(m1));
 endmodule

 module m_17 (
    input i1,
    input i2,
    input i3,
    input i4,
    output o1
 );
 wire m1;
 wire m2;
 wire m3;
 m_3 inst_1(.i1(m2),
           .o1(o1));
 m_11 inst_2(.i1(m3),
            .i2(m1),
            .o1(m2));
 m_9 inst_3(.i1(i3),
           .i2(i4),
           .o1(m1));
 m_9 inst_4(.i1(i1),
           .i2(i2),
           .o1(m3));
 endmodule

 module m_16 (
    input i1,
    input i2,
    output o1
 );
 m_9 inst_1(.i1(i1),
           .i2(i2),
           .o1(o1));
 endmodule

 module m_15 (
    input i1,
    input i2,
    output o1
 );
 m_11 inst_1(.i1(i1),
            .i2(i2),
            .o1(o1));
 endmodule

 module m_14 (
    input i1,
    input i2,
    input i3,
    output o1
 );
 wire m1;
 wire m2;
 m_3 inst_1(.i1(m1),
           .o1(o1));
 m_9 inst_2(.i1(m2),
           .i2(i3),
           .o1(m1));
 m_11 inst_3(.i1(i1),
            .i2(i2),
            .o1(m2));
 endmodule

 module m_13 (
    input i1,
    input i2,
    input i3,
    output o1
 );
 wire m1;
 wire m2;
 m_3 inst_1(.i1(m2),
           .o1(o1));
 m_11 inst_2(.i1(m1),
            .i2(i3),
            .o1(m2));
 m_11 inst_3(.i1(i1),
            .i2(i2),
            .o1(m1));
 endmodule

 module m_12 (
    input i1,
    input i2,
    input i3,
    output o1
 );
 wire m1;
 wire m2;
 m_3 inst_1(.i1(m1),
           .o1(o1));
 m_11 inst_2(.i1(m2),
            .i2(i3),
            .o1(m1));
 m_9 inst_3(.i1(i1),
           .i2(i2),
           .o1(m2));
 endmodule

 module m_10 (
    input i1,
    input i2,
    output o1
 );
 wire m1;
 m_3 inst_1(.i1(m1),
           .o1(o1));
 m_11 inst_2(.i1(i1),
            .i2(i2),
            .o1(m1));
 endmodule

 module m_11 (
    input i1,
    input i2,
    output o1
 );
 assign o1 = i1 & i2;
 endmodule

 module m_8 (
    input i1,
    input i2,
    output o1
 );
 wire m1;
 m_3 inst_1(.i1(m1),
           .o1(o1));
 m_9 inst_2(.i1(i1),
           .i2(i2),
           .o1(m1));
 endmodule

 module m_9 (
    input i1,
    input i2,
    output o1
 );
 assign o1 = i1 | i2;
 endmodule

 module m_6 (
    input i1,
    input i2,
    output o1
 );
 wire m1;
 m_3 inst_1(.i1(m1),
           .o1(o1));
 m_7 inst_2(.i1(i1),
           .i2(i2),
           .o1(m1));
 endmodule

 module m_7 (
    input i1,
    input i2,
    output o1
 );
 assign o1 = ~(i1) & i2 | i1 & ~(i2);
 endmodule

 module m_5 (
    input i1,
    output o1
 );
 m_3 inst_1(.i1(i1),
           .o1(o1));
 endmodule

 module m_2 (
    input i1,
    input i2,
    input i3,
    output o1
 );
 wire m1;
 m_4 inst_1(.i1(i3),
           .i2(i1),
           .i3(i2),
           .o1(m1));
 m_3 inst_2(.i1(m1),
           .o1(o1));
 endmodule

 module m_4 (
    input i1,
    input i2,
    input i3,
    output o1
 );
 assign o1 = i1 ? i2 : i3;
 endmodule

 module m_3 (
    input i1,
    output o1
 );
 assign o1 = ~(i1);
 endmodule

 module m_1 (
    input i1,
    output o1
 );
 assign o1 = i1;
 endmodule

 module m (
    input [1 : 0] i1,
    output [1 : 0] o1
 );
 assign o1 = i1[1:0];
 endmodule

