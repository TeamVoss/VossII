 module _synth_1 (
    input [1 : 0] i1,
    input i2,
    input [30 : 0] i3,
    input [30 : 0] i4,
    output [32 : 0] o1,
    output [8 : 0] o2,
    output o3,
    output [2 : 0] o4
 );
 wire m16;
 wire m1;
 wire m2;
 wire m3;
 wire m4;
 wire m5;
 wire [23 : 0] m6;
 wire [4 : 0] m7;
 wire [32 : 0] m8;
 wire [8 : 0] m9;
 wire [23 : 0] m10;
 wire [23 : 0] m11;
 wire [8 : 0] m12;
 wire [4 : 0] m13;
 wire [4 : 0] m14;
 wire [1 : 0] m15;
 m_9 inst_1(.i1(m5),
           .i2(m16),
           .o1(o3));
 m_8 inst_2(.i1(m12[7:5]),
           .o1(m16));
 m_8 inst_3(.i1(o2[7:5]),
           .o1(m1));
 m_8 inst_4(.i1(m9[7:5]),
           .o1(m2));
 m_7 inst_5(.i1(m11[7:0]),
           .o1(m3));
 m_6 inst_6(.i1(m8[8:0]),
           .o1(m4));
 m_5 inst_7(.i1(m12[8]),
           .o1(m5));
 m_4 inst_8(.i1(9'b010011101),
           .i2({1'b0, i3[30:23]}),
           .o1(m12[8:0]));
 m_4 inst_9(.i1({1'b0, i4[30:23]}),
           .i2({1'b0, i3[30:23]}),
           .o1(o2[8:0]));
 m_4 inst_10(.i1({1'b0, i3[30:23]}),
            .i2({1'b0, i4[30:23]}),
            .o1(m9[8:0]));
 m_2 inst_11(.i1(m1),
            .i2(5'b11111),
            .i3(o2[4:0]),
            .o1(m13[4:0]));
 m_2 inst_12(.i1(m2),
            .i2(5'b11111),
            .i3(m9[4:0]),
            .o1(m14[4:0]));
 m_3 inst_13(.i1(o2[8]),
            .i2({i1[1], i4[22:0]}),
            .i3({i1[0], i3[22:0]}),
            .o1(m10[23:0]));
 m_3 inst_14(.i1(o3),
            .i2(24'b000000000000000000000000),
            .i3({i1[0], i3[22:0]}),
            .o1(m6[23:0]));
 m_3 inst_15(.i1(i2),
            .i2(m6[23:0]),
            .i3(m10[23:0]),
            .o1(m11[23:0]));
 m_2 inst_16(.i1(o2[8]),
            .i2(m14[4:0]),
            .i3(m13[4:0]),
            .o1(m7[4:0]));
 m_2 inst_17(.i1(i2),
            .i2(m12[4:0]),
            .i3(m7[4:0]),
            .o1({m15[1:0], o4[2:0]}));
 m_1 inst_18(.i1(m15[1]),
            .i2({16'b0000000000000000, m11[23:8], m3}),
            .i3({m11[23:0], 9'b000000000}),
            .o1(m8[32:0]));
 m inst_19(.i1(m15[0]),
          .i2({8'b00000000, m8[32:9], m4}),
          .i3(m8[32:0]),
          .o1(o1[32:0]));
 endmodule

 module m_9 (
    input i1,
    input i2,
    output o1
 );
 assign o1 = i1 & i2;
 endmodule

 module m_8 (
    input [2 : 0] i1,
    output o1
 );
 assign o1 = ~(i1[2:0] == 3'b000);
 endmodule

 module m_7 (
    input [7 : 0] i1,
    output o1
 );
 assign o1 = ~(i1[7:0] == 8'b00000000);
 endmodule

 module m_6 (
    input [8 : 0] i1,
    output o1
 );
 assign o1 = ~(i1[8:0] == 9'b000000000);
 endmodule

 module m_5 (
    input i1,
    output o1
 );
 assign o1 = ~(i1);
 endmodule

 module m_4 (
    input [8 : 0] i1,
    input [8 : 0] i2,
    output [8 : 0] o1
 );
 assign o1 = i1[8:0] - i2[8:0];
 endmodule

 module m_3 (
    input i1,
    input [23 : 0] i2,
    input [23 : 0] i3,
    output [23 : 0] o1
 );
 assign o1 = i1 ? i2[23:0] : i3[23:0];
 endmodule

 module m_2 (
    input i1,
    input [4 : 0] i2,
    input [4 : 0] i3,
    output [4 : 0] o1
 );
 assign o1 = i1 ? i2[4:0] : i3[4:0];
 endmodule

 module m_1 (
    input i1,
    input [32 : 0] i2,
    input [32 : 0] i3,
    output [32 : 0] o1
 );
 assign o1 = i1 ? i2[32:0] : i3[32:0];
 endmodule

 module m (
    input i1,
    input [32 : 0] i2,
    input [32 : 0] i3,
    output [32 : 0] o1
 );
 assign o1 = i1 ? i2[32:0] : i3[32:0];
 endmodule

