 module _synth_103 (
    input i1,
    input [10 : 0] i2,
    input i3,
    input [30 : 0] i4,
    output [35 : 0] o1
 );
 wire [14 : 0] m2;
 wire m1;
 m_18 inst_1(.o1(m2[14:0]));
 m_17 inst_2(.o1(m1));
 mapped_adder inst_3(.i1(i1),
                    .i2({m2[14:0], i2[10:0]}),
                    .i3(i3),
                    .i4({i4[30:23], m1, i4[22:0]}),
                    .o1(o1[35:0]));
 endmodule

 module m_18 ( output [14 : 0] o1
 );
 assign o1 = 15'b000000000000000;
 endmodule

 module m_17 ( output o1
 );
 assign o1 = 1'b1;
 endmodule

 module mapped_adder (
    input i1,
    input [25 : 0] i2,
    input i3,
    input [31 : 0] i4,
    output [35 : 0] o1
 );
 wire m179;
 wire m1;
 wire m2;
 wire m3;
 wire m4;
 wire m5;
 wire m6;
 wire m7;
 wire m8;
 wire m9;
 wire m10;
 wire m11;
 wire m12;
 wire m13;
 wire m14;
 wire m15;
 wire m16;
 wire m17;
 wire m18;
 wire m19;
 wire m20;
 wire m21;
 wire m22;
 wire m23;
 wire m24;
 wire m25;
 wire m26;
 wire m27;
 wire m28;
 wire m29;
 wire m30;
 wire m31;
 wire m32;
 wire m33;
 wire m34;
 wire m35;
 wire m36;
 wire m37;
 wire m38;
 wire m39;
 wire m40;
 wire m41;
 wire m42;
 wire m43;
 wire m44;
 wire m45;
 wire m46;
 wire m47;
 wire m48;
 wire m49;
 wire m50;
 wire m51;
 wire m52;
 wire m53;
 wire m54;
 wire m55;
 wire m56;
 wire m57;
 wire m58;
 wire m59;
 wire m60;
 wire m61;
 wire m62;
 wire m63;
 wire m64;
 wire m65;
 wire m66;
 wire m67;
 wire m68;
 wire m69;
 wire m70;
 wire m71;
 wire m72;
 wire m73;
 wire m74;
 wire m75;
 wire m76;
 wire m77;
 wire m78;
 wire m79;
 wire m80;
 wire m81;
 wire m82;
 wire m83;
 wire m84;
 wire m85;
 wire m86;
 wire m87;
 wire m88;
 wire m89;
 wire m90;
 wire m91;
 wire m92;
 wire m93;
 wire m94;
 wire m95;
 wire m96;
 wire m97;
 wire m98;
 wire m99;
 wire m100;
 wire m101;
 wire m102;
 wire m103;
 wire m104;
 wire m105;
 wire m106;
 wire m107;
 wire m108;
 wire m109;
 wire m110;
 wire m111;
 wire m112;
 wire m113;
 wire m114;
 wire m115;
 wire m116;
 wire m117;
 wire m118;
 wire m119;
 wire m120;
 wire m121;
 wire m122;
 wire m123;
 wire m124;
 wire m125;
 wire m126;
 wire m127;
 wire m128;
 wire m129;
 wire m130;
 wire m131;
 wire m132;
 wire m133;
 wire m134;
 wire m135;
 wire m136;
 wire m137;
 wire m138;
 wire m139;
 wire m140;
 wire m141;
 wire m142;
 wire m143;
 wire m144;
 wire m145;
 wire m146;
 wire m147;
 wire m148;
 wire m149;
 wire m150;
 wire m151;
 wire m152;
 wire m153;
 wire m154;
 wire m155;
 wire m156;
 wire m157;
 wire m158;
 wire m159;
 wire m160;
 wire m161;
 wire m162;
 wire m163;
 wire m164;
 wire m165;
 wire m166;
 wire m167;
 wire m168;
 wire m169;
 wire m170;
 wire m171;
 wire m172;
 wire m173;
 wire m174;
 wire m175;
 wire m176;
 wire m177;
 wire m178;
 m_4 inst_1(.i1(i3),
           .o1(m179));
 m_15 inst_2(.i1(m179),
            .i2(m1),
            .i3(m2),
            .o1(o1[1]));
 m_10 inst_3(.i1(i1),
            .i2(i2[0]),
            .o1(m2));
 m_14 inst_4(.i1(m179),
            .i2(m3),
            .i3(m2),
            .o1(m4));
 m_4 inst_5(.i1(i2[1]),
           .o1(m3));
 m_5 inst_6(.i1(m4),
           .i2(m5),
           .i3(m7),
           .o1(m8));
 m_10 inst_7(.i1(i4[0]),
            .i2(m6),
            .o1(m5));
 m_1 inst_8(.i1(i1),
           .i2(i2[2]),
           .o1(m6));
 m_9 inst_9(.i1(i4[0]),
           .i2(m6),
           .o1(m7));
 m_5 inst_10(.i1(m9),
            .i2(m8),
            .i3(m10),
            .o1(m12));
 m_12 inst_11(.i1(i4[1]),
             .i2(m11),
             .o1(m9));
 m_13 inst_12(.i1(i4[1]),
             .i2(m11),
             .o1(m10));
 m_1 inst_13(.i1(i1),
            .i2(i2[3]),
            .o1(m11));
 m_5 inst_14(.i1(m13),
            .i2(m12),
            .i3(m15),
            .o1(m16));
 m_10 inst_15(.i1(i4[2]),
             .i2(m14),
             .o1(m13));
 m_1 inst_16(.i1(i1),
            .i2(i2[4]),
            .o1(m14));
 m_9 inst_17(.i1(i4[2]),
            .i2(m14),
            .o1(m15));
 m_5 inst_18(.i1(m17),
            .i2(m16),
            .i3(m18),
            .o1(m20));
 m_12 inst_19(.i1(i4[3]),
             .i2(m19),
             .o1(m17));
 m_13 inst_20(.i1(i4[3]),
             .i2(m19),
             .o1(m18));
 m_1 inst_21(.i1(i1),
            .i2(i2[5]),
            .o1(m19));
 m_5 inst_22(.i1(m21),
            .i2(m20),
            .i3(m23),
            .o1(m24));
 m_10 inst_23(.i1(i4[4]),
             .i2(m22),
             .o1(m21));
 m_1 inst_24(.i1(i1),
            .i2(i2[6]),
            .o1(m22));
 m_9 inst_25(.i1(i4[4]),
            .i2(m22),
            .o1(m23));
 m_5 inst_26(.i1(m25),
            .i2(m24),
            .i3(m26),
            .o1(m28));
 m_12 inst_27(.i1(i4[5]),
             .i2(m27),
             .o1(m25));
 m_13 inst_28(.i1(i4[5]),
             .i2(m27),
             .o1(m26));
 m_1 inst_29(.i1(i1),
            .i2(i2[7]),
            .o1(m27));
 m_5 inst_30(.i1(m29),
            .i2(m28),
            .i3(m31),
            .o1(m32));
 m_10 inst_31(.i1(i4[6]),
             .i2(m30),
             .o1(m29));
 m_1 inst_32(.i1(i1),
            .i2(i2[8]),
            .o1(m30));
 m_9 inst_33(.i1(i4[6]),
            .i2(m30),
            .o1(m31));
 m_5 inst_34(.i1(m33),
            .i2(m32),
            .i3(m34),
            .o1(m36));
 m_12 inst_35(.i1(i4[7]),
             .i2(m35),
             .o1(m33));
 m_13 inst_36(.i1(i4[7]),
             .i2(m35),
             .o1(m34));
 m_1 inst_37(.i1(i1),
            .i2(i2[9]),
            .o1(m35));
 m_5 inst_38(.i1(m37),
            .i2(m36),
            .i3(m39),
            .o1(m40));
 m_10 inst_39(.i1(i4[8]),
             .i2(m38),
             .o1(m37));
 m_1 inst_40(.i1(i1),
            .i2(i2[10]),
            .o1(m38));
 m_9 inst_41(.i1(i4[8]),
            .i2(m38),
            .o1(m39));
 m_5 inst_42(.i1(m41),
            .i2(m40),
            .i3(m42),
            .o1(m44));
 m_12 inst_43(.i1(i4[9]),
             .i2(m43),
             .o1(m41));
 m_13 inst_44(.i1(i4[9]),
             .i2(m43),
             .o1(m42));
 m_1 inst_45(.i1(i1),
            .i2(i2[11]),
            .o1(m43));
 m_11 inst_46(.i1(m45),
             .i2(m44),
             .i3(m46),
             .o1(m48));
 m_9 inst_47(.i1(i4[10]),
            .i2(m47),
            .o1(m45));
 m_10 inst_48(.i1(i4[10]),
             .i2(m47),
             .o1(m46));
 m_1 inst_49(.i1(i1),
            .i2(i2[12]),
            .o1(m47));
 m_5 inst_50(.i1(m49),
            .i2(m48),
            .i3(m50),
            .o1(m52));
 m_12 inst_51(.i1(i4[11]),
             .i2(m51),
             .o1(m49));
 m_13 inst_52(.i1(i4[11]),
             .i2(m51),
             .o1(m50));
 m_1 inst_53(.i1(i1),
            .i2(i2[13]),
            .o1(m51));
 m_11 inst_54(.i1(m53),
             .i2(m52),
             .i3(m54),
             .o1(m56));
 m_9 inst_55(.i1(i4[12]),
            .i2(m55),
            .o1(m53));
 m_10 inst_56(.i1(i4[12]),
             .i2(m55),
             .o1(m54));
 m_1 inst_57(.i1(i1),
            .i2(i2[14]),
            .o1(m55));
 m_11 inst_58(.i1(m57),
             .i2(m56),
             .i3(m59),
             .o1(m60));
 m_13 inst_59(.i1(i4[13]),
             .i2(m58),
             .o1(m57));
 m_1 inst_60(.i1(i1),
            .i2(i2[15]),
            .o1(m58));
 m_12 inst_61(.i1(i4[13]),
             .i2(m58),
             .o1(m59));
 m_5 inst_62(.i1(m61),
            .i2(m60),
            .i3(m63),
            .o1(m64));
 m_10 inst_63(.i1(i4[14]),
             .i2(m62),
             .o1(m61));
 m_1 inst_64(.i1(i1),
            .i2(i2[16]),
            .o1(m62));
 m_9 inst_65(.i1(i4[14]),
            .i2(m62),
            .o1(m63));
 m_11 inst_66(.i1(m65),
             .i2(m64),
             .i3(m67),
             .o1(m68));
 m_13 inst_67(.i1(i4[15]),
             .i2(m66),
             .o1(m65));
 m_1 inst_68(.i1(i1),
            .i2(i2[17]),
            .o1(m66));
 m_12 inst_69(.i1(i4[15]),
             .i2(m66),
             .o1(m67));
 m_5 inst_70(.i1(m69),
            .i2(m68),
            .i3(m71),
            .o1(m72));
 m_10 inst_71(.i1(i4[16]),
             .i2(m70),
             .o1(m69));
 m_1 inst_72(.i1(i1),
            .i2(i2[18]),
            .o1(m70));
 m_9 inst_73(.i1(i4[16]),
            .i2(m70),
            .o1(m71));
 m_11 inst_74(.i1(m73),
             .i2(m72),
             .i3(m75),
             .o1(m76));
 m_13 inst_75(.i1(i4[17]),
             .i2(m74),
             .o1(m73));
 m_1 inst_76(.i1(i1),
            .i2(i2[19]),
            .o1(m74));
 m_12 inst_77(.i1(i4[17]),
             .i2(m74),
             .o1(m75));
 m_5 inst_78(.i1(m77),
            .i2(m76),
            .i3(m79),
            .o1(m80));
 m_10 inst_79(.i1(i4[18]),
             .i2(m78),
             .o1(m77));
 m_1 inst_80(.i1(i1),
            .i2(i2[20]),
            .o1(m78));
 m_9 inst_81(.i1(i4[18]),
            .i2(m78),
            .o1(m79));
 m_11 inst_82(.i1(m81),
             .i2(m80),
             .i3(m83),
             .o1(m84));
 m_13 inst_83(.i1(i4[19]),
             .i2(m82),
             .o1(m81));
 m_1 inst_84(.i1(i1),
            .i2(i2[21]),
            .o1(m82));
 m_12 inst_85(.i1(i4[19]),
             .i2(m82),
             .o1(m83));
 m_5 inst_86(.i1(m85),
            .i2(m84),
            .i3(m87),
            .o1(m88));
 m_10 inst_87(.i1(i4[20]),
             .i2(m86),
             .o1(m85));
 m_1 inst_88(.i1(i1),
            .i2(i2[22]),
            .o1(m86));
 m_9 inst_89(.i1(i4[20]),
            .i2(m86),
            .o1(m87));
 m_11 inst_90(.i1(m89),
             .i2(m88),
             .i3(m91),
             .o1(m92));
 m_13 inst_91(.i1(i4[21]),
             .i2(m90),
             .o1(m89));
 m_1 inst_92(.i1(i1),
            .i2(i2[23]),
            .o1(m90));
 m_12 inst_93(.i1(i4[21]),
             .i2(m90),
             .o1(m91));
 m_5 inst_94(.i1(m93),
            .i2(m92),
            .i3(m95),
            .o1(m96));
 m_10 inst_95(.i1(i4[22]),
             .i2(m94),
             .o1(m93));
 m_1 inst_96(.i1(i1),
            .i2(i2[24]),
            .o1(m94));
 m_9 inst_97(.i1(i4[22]),
            .i2(m94),
            .o1(m95));
 m_11 inst_98(.i1(m97),
             .i2(m96),
             .i3(m99),
             .o1(m100));
 m_13 inst_99(.i1(i4[23]),
             .i2(m98),
             .o1(m97));
 m_1 inst_100(.i1(i1),
             .i2(i2[25]),
             .o1(m98));
 m_12 inst_101(.i1(i4[23]),
              .i2(m98),
              .o1(m99));
 m_5 inst_102(.i1(m101),
             .i2(m100),
             .i3(m102),
             .o1(m103));
 m_10 inst_103(.i1(m177),
              .i2(i4[24]),
              .o1(m101));
 m_9 inst_104(.i1(m177),
             .i2(i4[24]),
             .o1(m102));
 m_11 inst_105(.i1(m104),
              .i2(m103),
              .i3(m105),
              .o1(m107));
 m_9 inst_106(.i1(i1),
             .i2(m106),
             .o1(m104));
 m_10 inst_107(.i1(i1),
              .i2(m106),
              .o1(m105));
 m_4 inst_108(.i1(i4[25]),
             .o1(m106));
 m_11 inst_109(.i1(m108),
              .i2(m107),
              .i3(m109),
              .o1(m110));
 m_9 inst_110(.i1(m177),
             .i2(i4[26]),
             .o1(m108));
 m_10 inst_111(.i1(m177),
              .i2(i4[26]),
              .o1(m109));
 m_5 inst_112(.i1(m111),
             .i2(m110),
             .i3(m113),
             .o1(m114));
 m_10 inst_113(.i1(i1),
              .i2(m112),
              .o1(m111));
 m_4 inst_114(.i1(i4[27]),
             .o1(m112));
 m_9 inst_115(.i1(i1),
             .i2(m112),
             .o1(m113));
 m_5 inst_116(.i1(m115),
             .i2(m114),
             .i3(m116),
             .o1(m117));
 m_10 inst_117(.i1(m177),
              .i2(i4[28]),
              .o1(m115));
 m_9 inst_118(.i1(m177),
             .i2(i4[28]),
             .o1(m116));
 m_11 inst_119(.i1(m118),
              .i2(m117),
              .i3(m119),
              .o1(m121));
 m_9 inst_120(.i1(i1),
             .i2(m120),
             .o1(m118));
 m_10 inst_121(.i1(i1),
              .i2(m120),
              .o1(m119));
 m_4 inst_122(.i1(i4[29]),
             .o1(m120));
 m_5 inst_123(.i1(m126),
             .i2(m121),
             .i3(i1),
             .o1(m128));
 m_5 inst_124(.i1(m122),
             .i2(m121),
             .i3(m123),
             .o1(m124));
 m_10 inst_125(.i1(m177),
              .i2(i4[30]),
              .o1(m122));
 m_9 inst_126(.i1(m177),
             .i2(i4[30]),
             .o1(m123));
 m_11 inst_127(.i1(m129),
              .i2(m124),
              .i3(m130),
              .o1(o1[35]));
 m_1 inst_128(.i1(m124),
             .i2(m125),
             .o1(o1[34]));
 m_8 inst_129(.i1(i1),
             .i2(i4[31]),
             .o1(m125));
 m_4 inst_130(.i1(i4[30]),
             .o1(m126));
 m_10 inst_131(.i1(i1),
              .i2(m126),
              .o1(m127));
 m_5 inst_132(.i1(i1),
             .i2(m129),
             .i3(m128),
             .o1(m130));
 m_4 inst_133(.i1(i4[31]),
             .o1(m129));
 m_1 inst_134(.i1(m121),
             .i2(m131),
             .o1(o1[33]));
 m_10 inst_135(.i1(m122),
              .i2(m127),
              .o1(m131));
 m_1 inst_136(.i1(m132),
             .i2(m117),
             .o1(o1[32]));
 m_9 inst_137(.i1(m133),
             .i2(m118),
             .o1(m132));
 m_9 inst_138(.i1(m177),
             .i2(i4[29]),
             .o1(m133));
 m_1 inst_139(.i1(m114),
             .i2(m134),
             .o1(o1[31]));
 m_1 inst_140(.i1(i1),
             .i2(i4[28]),
             .o1(m134));
 m_1 inst_141(.i1(m110),
             .i2(m135),
             .o1(o1[30]));
 m_9 inst_142(.i1(m136),
             .i2(m113),
             .o1(m135));
 m_9 inst_143(.i1(m177),
             .i2(i4[27]),
             .o1(m136));
 m_1 inst_144(.i1(m107),
             .i2(m137),
             .o1(o1[29]));
 m_1 inst_145(.i1(i1),
             .i2(i4[26]),
             .o1(m137));
 m_1 inst_146(.i1(m138),
             .i2(m103),
             .o1(o1[28]));
 m_9 inst_147(.i1(m139),
             .i2(m104),
             .o1(m138));
 m_9 inst_148(.i1(m177),
             .i2(i4[25]),
             .o1(m139));
 m_1 inst_149(.i1(m100),
             .i2(m140),
             .o1(o1[27]));
 m_1 inst_150(.i1(i1),
             .i2(i4[24]),
             .o1(m140));
 m_1 inst_151(.i1(m141),
             .i2(m96),
             .o1(o1[26]));
 m_9 inst_152(.i1(m142),
             .i2(m97),
             .o1(m141));
 m_9 inst_153(.i1(i4[23]),
             .i2(m98),
             .o1(m142));
 m_1 inst_154(.i1(m92),
             .i2(m143),
             .o1(o1[25]));
 m_8 inst_155(.i1(i4[22]),
             .i2(m94),
             .o1(m143));
 m_1 inst_156(.i1(m144),
             .i2(m88),
             .o1(o1[24]));
 m_9 inst_157(.i1(m145),
             .i2(m89),
             .o1(m144));
 m_9 inst_158(.i1(i4[21]),
             .i2(m90),
             .o1(m145));
 m_1 inst_159(.i1(m84),
             .i2(m146),
             .o1(o1[23]));
 m_8 inst_160(.i1(i4[20]),
             .i2(m86),
             .o1(m146));
 m_1 inst_161(.i1(m147),
             .i2(m80),
             .o1(o1[22]));
 m_9 inst_162(.i1(m81),
             .i2(m148),
             .o1(m147));
 m_9 inst_163(.i1(i4[19]),
             .i2(m82),
             .o1(m148));
 m_1 inst_164(.i1(m76),
             .i2(m149),
             .o1(o1[21]));
 m_8 inst_165(.i1(i4[18]),
             .i2(m78),
             .o1(m149));
 m_1 inst_166(.i1(m150),
             .i2(m72),
             .o1(o1[20]));
 m_9 inst_167(.i1(m151),
             .i2(m73),
             .o1(m150));
 m_9 inst_168(.i1(i4[17]),
             .i2(m74),
             .o1(m151));
 m_1 inst_169(.i1(m68),
             .i2(m152),
             .o1(o1[19]));
 m_8 inst_170(.i1(i4[16]),
             .i2(m70),
             .o1(m152));
 m_1 inst_171(.i1(m153),
             .i2(m64),
             .o1(o1[18]));
 m_9 inst_172(.i1(m154),
             .i2(m65),
             .o1(m153));
 m_9 inst_173(.i1(i4[15]),
             .i2(m66),
             .o1(m154));
 m_1 inst_174(.i1(m60),
             .i2(m155),
             .o1(o1[17]));
 m_8 inst_175(.i1(i4[14]),
             .i2(m62),
             .o1(m155));
 m_1 inst_176(.i1(m156),
             .i2(m56),
             .o1(o1[16]));
 m_9 inst_177(.i1(m157),
             .i2(m57),
             .o1(m156));
 m_9 inst_178(.i1(i4[13]),
             .i2(m58),
             .o1(m157));
 m_1 inst_179(.i1(m52),
             .i2(m158),
             .o1(o1[15]));
 m_8 inst_180(.i1(i4[12]),
             .i2(m55),
             .o1(m158));
 m_1 inst_181(.i1(m48),
             .i2(m159),
             .o1(o1[14]));
 m_9 inst_182(.i1(m160),
             .i2(m50),
             .o1(m159));
 m_9 inst_183(.i1(i4[11]),
             .i2(m51),
             .o1(m160));
 m_1 inst_184(.i1(m44),
             .i2(m161),
             .o1(o1[13]));
 m_8 inst_185(.i1(i4[10]),
             .i2(m47),
             .o1(m161));
 m_1 inst_186(.i1(m40),
             .i2(m162),
             .o1(o1[12]));
 m_9 inst_187(.i1(m163),
             .i2(m42),
             .o1(m162));
 m_9 inst_188(.i1(i4[9]),
             .i2(m43),
             .o1(m163));
 m_1 inst_189(.i1(m164),
             .i2(m36),
             .o1(o1[11]));
 m_8 inst_190(.i1(i4[8]),
             .i2(m38),
             .o1(m164));
 m_1 inst_191(.i1(m32),
             .i2(m165),
             .o1(o1[10]));
 m_9 inst_192(.i1(m166),
             .i2(m34),
             .o1(m165));
 m_9 inst_193(.i1(i4[7]),
             .i2(m35),
             .o1(m166));
 m_1 inst_194(.i1(m167),
             .i2(m28),
             .o1(o1[9]));
 m_8 inst_195(.i1(i4[6]),
             .i2(m30),
             .o1(m167));
 m_1 inst_196(.i1(m24),
             .i2(m168),
             .o1(o1[8]));
 m_9 inst_197(.i1(m169),
             .i2(m26),
             .o1(m168));
 m_9 inst_198(.i1(i4[5]),
             .i2(m27),
             .o1(m169));
 m_1 inst_199(.i1(m170),
             .i2(m20),
             .o1(o1[7]));
 m_8 inst_200(.i1(i4[4]),
             .i2(m22),
             .o1(m170));
 m_1 inst_201(.i1(m16),
             .i2(m171),
             .o1(o1[6]));
 m_9 inst_202(.i1(m172),
             .i2(m18),
             .o1(m171));
 m_9 inst_203(.i1(i4[3]),
             .i2(m19),
             .o1(m172));
 m_1 inst_204(.i1(m173),
             .i2(m12),
             .o1(o1[5]));
 m_8 inst_205(.i1(i4[2]),
             .i2(m14),
             .o1(m173));
 m_1 inst_206(.i1(m8),
             .i2(m174),
             .o1(o1[4]));
 m_9 inst_207(.i1(m175),
             .i2(m10),
             .o1(m174));
 m_9 inst_208(.i1(i4[1]),
             .i2(m11),
             .o1(m175));
 m_1 inst_209(.i1(m4),
             .i2(m176),
             .o1(o1[3]));
 m_8 inst_210(.i1(i4[0]),
             .i2(m6),
             .o1(m176));
 m_5 inst_211(.i1(i1),
             .i2(m179),
             .i3(i2[0]),
             .o1(m1));
 m_5 inst_212(.i1(i3),
             .i2(i2[0]),
             .i3(m177),
             .o1(m178));
 m_4 inst_213(.i1(i1),
             .o1(m177));
 m_1 inst_214(.i1(i2[1]),
             .i2(m178),
             .o1(o1[2]));
 m inst_215(.i1(i3),
           .o1(o1[0]));
 endmodule

 module m_15 (
    input i1,
    input i2,
    input i3,
    output o1
 );
 wire m1;
 m_16 inst_1(.i1(i3),
            .i2(i1),
            .i3(i2),
            .o1(m1));
 m_3 inst_2(.i1(m1),
           .o1(o1));
 endmodule

 module m_16 (
    input i1,
    input i2,
    input i3,
    output o1
 );
 assign o1 = i1 ? i2 : i3;
 endmodule

 module m_14 (
    input i1,
    input i2,
    input i3,
    output o1
 );
 wire m1;
 wire m2;
 m_3 inst_1(.i1(m2),
           .o1(o1));
 m_7 inst_2(.i1(m1),
           .i2(i3),
           .o1(m2));
 m_7 inst_3(.i1(i1),
           .i2(i2),
           .o1(m1));
 endmodule

 module m_13 (
    input i1,
    input i2,
    output o1
 );
 m_6 inst_1(.i1(i1),
           .i2(i2),
           .o1(o1));
 endmodule

 module m_12 (
    input i1,
    input i2,
    output o1
 );
 m_7 inst_1(.i1(i1),
           .i2(i2),
           .o1(o1));
 endmodule

 module m_11 (
    input i1,
    input i2,
    input i3,
    output o1
 );
 wire m1;
 wire m2;
 m_3 inst_1(.i1(m1),
           .o1(o1));
 m_6 inst_2(.i1(m2),
           .i2(i3),
           .o1(m1));
 m_7 inst_3(.i1(i1),
           .i2(i2),
           .o1(m2));
 endmodule

 module m_10 (
    input i1,
    input i2,
    output o1
 );
 wire m1;
 m_3 inst_1(.i1(m1),
           .o1(o1));
 m_6 inst_2(.i1(i1),
           .i2(i2),
           .o1(m1));
 endmodule

 module m_9 (
    input i1,
    input i2,
    output o1
 );
 wire m1;
 m_3 inst_1(.i1(m1),
           .o1(o1));
 m_7 inst_2(.i1(i1),
           .i2(i2),
           .o1(m1));
 endmodule

 module m_8 (
    input i1,
    input i2,
    output o1
 );
 m_2 inst_1(.i1(i1),
           .i2(i2),
           .o1(o1));
 endmodule

 module m_5 (
    input i1,
    input i2,
    input i3,
    output o1
 );
 wire m1;
 wire m2;
 m_3 inst_1(.i1(m1),
           .o1(o1));
 m_7 inst_2(.i1(m2),
           .i2(i3),
           .o1(m1));
 m_6 inst_3(.i1(i1),
           .i2(i2),
           .o1(m2));
 endmodule

 module m_7 (
    input i1,
    input i2,
    output o1
 );
 assign o1 = i1 & i2;
 endmodule

 module m_6 (
    input i1,
    input i2,
    output o1
 );
 assign o1 = i1 | i2;
 endmodule

 module m_4 (
    input i1,
    output o1
 );
 m_3 inst_1(.i1(i1),
           .o1(o1));
 endmodule

 module m_1 (
    input i1,
    input i2,
    output o1
 );
 wire m1;
 m_3 inst_1(.i1(m1),
           .o1(o1));
 m_2 inst_2(.i1(i1),
           .i2(i2),
           .o1(m1));
 endmodule

 module m_3 (
    input i1,
    output o1
 );
 assign o1 = ~(i1);
 endmodule

 module m_2 (
    input i1,
    input i2,
    output o1
 );
 assign o1 = ~(i1) & i2 | i1 & ~(i2);
 endmodule

 module m (
    input i1,
    output o1
 );
 assign o1 = i1;
 endmodule

