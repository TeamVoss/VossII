 module _synth_31 (
    input [1 : 0] i1,
    input [1 : 0] i2,
    input [3 : 0] i3,
    input [31 : 0] i4,
    input [31 : 0] i5,
    input [33 : 0] i6,
    input [31 : 0] i7,
    input [36 : 0] i8,
    input [1 : 0] i9,
    input [35 : 0] i10,
    input [35 : 0] i11,
    input [1 : 0] i12,
    input i13,
    input i14,
    input [9 : 0] i15,
    input i16,
    input i17,
    input [35 : 0] i18,
    input i19,
    output [36 : 0] o1,
    output o2,
    output [31 : 0] o3,
    output [33 : 0] o4,
    output [31 : 0] o5,
    output [36 : 0] o6,
    output o7,
    output o8,
    output [9 : 0] o9,
    output o10,
    output o11,
    output o12,
    output o13,
    output [27 : 0] o14,
    output o15,
    output o16,
    output [31 : 0] o17,
    output o18,
    output o19,
    output [24 : 0] o20,
    output [24 : 0] o21
 );
 wire m126;
 wire m1;
 wire m2;
 wire m3;
 wire m4;
 wire m5;
 wire m6;
 wire m7;
 wire m8;
 wire m9;
 wire m10;
 wire m11;
 wire m12;
 wire m13;
 wire m14;
 wire m15;
 wire m16;
 wire m17;
 wire m18;
 wire m19;
 wire m20;
 wire m21;
 wire m22;
 wire m23;
 wire m24;
 wire m25;
 wire m26;
 wire m27;
 wire m28;
 wire m29;
 wire m30;
 wire m31;
 wire m32;
 wire m33;
 wire m34;
 wire m35;
 wire m36;
 wire m37;
 wire m38;
 wire m39;
 wire m40;
 wire m41;
 wire m42;
 wire m43;
 wire m44;
 wire m45;
 wire m46;
 wire m47;
 wire m48;
 wire m49;
 wire m50;
 wire m51;
 wire m52;
 wire m53;
 wire m54;
 wire m55;
 wire m56;
 wire m57;
 wire m58;
 wire m59;
 wire m60;
 wire m61;
 wire m62;
 wire [30 : 0] m63;
 wire m64;
 wire m65;
 wire m66;
 wire m67;
 wire m68;
 wire m69;
 wire m70;
 wire m71;
 wire m72;
 wire m73;
 wire m74;
 wire [9 : 0] m75;
 wire m76;
 wire [23 : 0] m77;
 wire [4 : 0] m78;
 wire m79;
 wire [32 : 0] m80;
 wire [31 : 0] m84;
 wire m81;
 wire m82;
 wire m83;
 wire [31 : 0] m85;
 wire [31 : 0] m86;
 wire [31 : 0] m87;
 wire [31 : 0] m88;
 wire [31 : 0] m89;
 wire [32 : 0] m90;
 wire [32 : 0] m91;
 wire [32 : 0] m92;
 wire [32 : 0] m93;
 wire [4 : 0] m94;
 wire m95;
 wire [7 : 0] m96;
 wire [8 : 0] m97;
 wire [8 : 0] m98;
 wire [9 : 0] m99;
 wire m100;
 wire [32 : 0] m101;
 wire [1 : 0] m102;
 wire [23 : 0] m103;
 wire m104;
 wire [31 : 0] m105;
 wire [31 : 0] m106;
 wire [23 : 0] m107;
 wire [36 : 0] m108;
 wire m109;
 wire m110;
 wire [23 : 0] m111;
 wire [35 : 0] m112;
 wire [8 : 0] m113;
 wire [8 : 0] m114;
 wire [4 : 0] m115;
 wire [4 : 0] m116;
 wire [4 : 0] m117;
 wire m118;
 wire m119;
 wire m120;
 wire m121;
 wire [33 : 0] m122;
 wire m123;
 wire [33 : 0] m124;
 wire m125;
 m_53 inst_1(.i1(m80[32:0]),
            .i2({32'b00000000000000000000000000000000, m95}),
            .o1(m101[32:0]));
 m_52 inst_2(.i1(m84[31:0]),
            .i2({31'b0000000000000000000000000000000, m105[31]}),
            .o1(m106[31:0]));
 m_51 inst_3(.i1(m64),
            .i2(m12),
            .o1(m1));
 m_51 inst_4(.i1(m1),
            .i2(m46),
            .o1(o7));
 m_51 inst_5(.i1(m47),
            .i2(m24),
            .o1(m100));
 m_51 inst_6(.i1(m49),
            .i2(m25),
            .o1(m2));
 m_51 inst_7(.i1(m50),
            .i2(m26),
            .o1(m3));
 m_51 inst_8(.i1(m51),
            .i2(m27),
            .o1(m4));
 m_51 inst_9(.i1(m13),
            .i2(i1[1]),
            .o1(m104));
 m_51 inst_10(.i1(m16),
             .i2(m103[23]),
             .o1(m5));
 m_51 inst_11(.i1(m52),
             .i2(m53),
             .o1(m6));
 m_51 inst_12(.i1(m54),
             .i2(m76),
             .o1(o2));
 m_51 inst_13(.i1(m56),
             .i2(m57),
             .o1(m7));
 m_51 inst_14(.i1(m7),
             .i2(m58),
             .o1(m8));
 m_51 inst_15(.i1(m59),
             .i2(m60),
             .o1(m9));
 m_51 inst_16(.i1(m19),
             .i2(m66),
             .o1(m10));
 m_51 inst_17(.i1(o13),
             .i2(m61),
             .o1(o8));
 m_51 inst_18(.i1(m62),
             .i2(m23),
             .o1(m11));
 m_41 inst_19(.i1(i3[1:0]),
             .o1(m12));
 m_50 inst_20(.i1(i4[31:0]),
             .o1(m13));
 m_46 inst_21(.i1(m98[8:1]),
             .o1(m14));
 m_49 inst_22(.i1(m98[8:0]),
             .o1(m15));
 m_46 inst_23(.i1(m98[7:0]),
             .o1(m16));
 m_48 inst_24(.i1(i4[31:0]),
             .i2(i5[31:0]),
             .o1(m17));
 m_47 inst_25(.i1(m85[31:16]),
             .o1(o19));
 m_46 inst_26(.i1(m86[31:24]),
             .o1(o18));
 m_45 inst_27(.i1(i7[31:28]),
             .o1(m120));
 m_24 inst_28(.i1(m87[31:30]),
             .o1(m119));
 m_41 inst_29(.i1(i3[1:0]),
             .o1(m18));
 m_44 inst_30(.i1(m85[31:0]),
             .o1(m19));
 m_43 inst_31(.i1(i3[1:0]),
             .o1(m20));
 m_42 inst_32(.i1({m94[0], o14[1:0]}),
             .o1(m21));
 m_41 inst_33(.i1(o14[1:0]),
             .o1(m22));
 m_24 inst_34(.i1(o14[1:0]),
             .o1(m23));
 m_40 inst_35(.i1(i18[26:0]),
             .o1(m125));
 m_33 inst_36(.i1(m113[7:5]),
             .o1(m24));
 m_36 inst_37(.i1(m114[7:3]),
             .o1(m25));
 m_39 inst_38(.i1(m114[7:4]),
             .o1(m26));
 m_33 inst_39(.i1(m114[7:5]),
             .o1(m27));
 m_34 inst_40(.i1(o17[24]),
             .i2(m112[27]),
             .o1(m28));
 m_33 inst_41(.i1(m112[2:0]),
             .o1(m29));
 m_32 inst_42(.i1(m112[1:0]),
             .o1(m30));
 m_35 inst_43(.i1(m89[6:0]),
             .o1(m31));
 m_33 inst_44(.i1(m98[7:5]),
             .o1(m32));
 m_33 inst_45(.i1(m97[7:5]),
             .o1(m33));
 m_38 inst_46(.i1(m111[7:0]),
             .o1(m34));
 m_37 inst_47(.i1(m90[8:0]),
             .o1(m35));
 m_36 inst_48(.i1(m91[4:0]),
             .o1(m36));
 m_33 inst_49(.i1(m92[2:0]),
             .o1(m37));
 m_32 inst_50(.i1(m93[1:0]),
             .o1(m38));
 m_34 inst_51(.i1(m101[8]),
             .i2(m101[7]),
             .o1(m39));
 m_34 inst_52(.i1(m101[16]),
             .i2(m101[15]),
             .o1(m40));
 m_34 inst_53(.i1(m101[32]),
             .i2(m101[31]),
             .o1(m41));
 m_35 inst_54(.i1({m94[4:0], o14[1:0]}),
             .o1(o16));
 m_34 inst_55(.i1(o17[24]),
             .i2(i18[27]),
             .o1(m42));
 m_33 inst_56(.i1(i18[2:0]),
             .o1(m43));
 m_32 inst_57(.i1(i18[1:0]),
             .o1(m44));
 m_32 inst_58(.i1(i18[1:0]),
             .o1(m45));
 m_31 inst_59(.i1(m104),
             .o1(m46));
 m_31 inst_60(.i1(m113[8]),
             .o1(m47));
 m_31 inst_61(.i1(i1[1]),
             .o1(m48));
 m_31 inst_62(.i1(m114[8]),
             .o1(m49));
 m_31 inst_63(.i1(m114[8]),
             .o1(m50));
 m_31 inst_64(.i1(m114[8]),
             .o1(m51));
 m_31 inst_65(.i1(m59),
             .o1(o13));
 m_31 inst_66(.i1(i2[1]),
             .o1(m52));
 m_31 inst_67(.i1(i2[0]),
             .o1(m53));
 m_31 inst_68(.i1(o15),
             .o1(m54));
 m_31 inst_69(.i1(i4[31]),
             .o1(m55));
 m_31 inst_70(.i1(m88[31]),
             .o1(m118));
 m_31 inst_71(.i1(i3[1]),
             .o1(m56));
 m_31 inst_72(.i1(i2[1]),
             .o1(m57));
 m_31 inst_73(.i1(i2[0]),
             .o1(m58));
 m_31 inst_74(.i1(i3[1]),
             .o1(m60));
 m_31 inst_75(.i1(i3[1]),
             .o1(m61));
 m_31 inst_76(.i1(m100),
             .o1(m62));
 m_30 inst_77(.i1({o14[27:2], m94[4:0]}),
             .o1(m63[30:0]));
 m_28 inst_78(.i1(m109),
             .i2(m110),
             .o1(m64));
 m_28 inst_79(.i1(m14),
             .i2(m15),
             .o1(m65));
 m_28 inst_80(.i1(m65),
             .i2(i3[1]),
             .o1(o11));
 m_28 inst_81(.i1(m98[8]),
             .i2(m5),
             .o1(m121));
 m_28 inst_82(.i1(m17),
             .i2(m6),
             .o1(o15));
 m_29 inst_83(.i1(m75[9:0]),
             .i2({1'b0, i13, 8'b00000000}),
             .o1(m99[9:0]));
 m_28 inst_84(.i1(m8),
             .i2(m10),
             .o1(o12));
 m_28 inst_85(.i1(m9),
             .i2(m20),
             .o1(m66));
 m_28 inst_86(.i1(m21),
             .i2(m22),
             .o1(m67));
 m_27 inst_87(.i1(m69),
             .i2(m39),
             .i3(m68),
             .i4(m40),
             .i5(m41),
             .o1(m110));
 m_25 inst_88(.i1(i1[1:0]),
             .o1(m68));
 m_24 inst_89(.i1(i1[1:0]),
             .o1(m69));
 m_27 inst_90(.i1(m70),
             .i2(m83),
             .i3(i3[3]),
             .i4(m79),
             .i5(i4[31]),
             .o1(m95));
 m_24 inst_91(.i1(i3[3:2]),
             .o1(m70));
 m_27 inst_92(.i1(m72),
             .i2(m2),
             .i3(m71),
             .i4(m3),
             .i5(m4),
             .o1(m109));
 m_25 inst_93(.i1(i1[1:0]),
             .o1(m71));
 m_24 inst_94(.i1(i1[1:0]),
             .o1(m72));
 m_26 inst_95(.i1(m74),
             .i2({i4[7], i4[7], i4[7], i4[7], i4[7], i4[7], i4[7], i4[7], i4[7], i4[7], i4[7], i4[7], i4[7], i4[7], i4[7], i4[7], i4[7], i4[7], i4[7], i4[7], i4[7], i4[7], i4[7], i4[7], i4[7:0]}),
             .i3(m73),
             .i4({i4[15], i4[15], i4[15], i4[15], i4[15], i4[15], i4[15], i4[15], i4[15], i4[15], i4[15], i4[15], i4[15], i4[15], i4[15], i4[15], i4[15:0]}),
             .i5(i4[31:0]),
             .o1(m105[31:0]));
 m_25 inst_96(.i1(i1[1:0]),
             .o1(m73));
 m_24 inst_97(.i1(i1[1:0]),
             .o1(m74));
 m_21 inst_98(.i1(9'b010011101),
             .i2({1'b0, i4[30:23]}),
             .o1(m113[8:0]));
 m_21 inst_99(.i1({1'b0, i4[30:23]}),
             .i2({8'b00111111, m48}),
             .o1(m114[8:0]));
 m_21 inst_100(.i1({1'b0, i5[30:23]}),
              .i2({1'b0, i4[30:23]}),
              .o1(m98[8:0]));
 m_23 inst_101(.i1({1'b0, i5[22:0]}),
              .i2({1'b0, i4[22:0]}),
              .o1(m103[23:0]));
 m_22 inst_102(.i1(i15[9:0]),
              .i2({5'b00000, i9[1:0], m120, m119, m118}),
              .o1(m75[9:0]));
 m_21 inst_103(.i1({1'b0, i4[30:23]}),
              .i2({1'b0, i5[30:23]}),
              .o1(m97[8:0]));
 m_20 inst_104(.i1(o17[31:24]),
              .i2(8'b00000001),
              .o1(m96[7:0]));
 m_19 inst_105(.i1(m98[0]),
              .i2({1'b0, i2[0], i4[22:0]}),
              .i3({i2[0], i4[22:0], 1'b0}),
              .o1(o20[24:0]));
 m_19 inst_106(.i1(m98[0]),
              .i2({1'b0, i2[1], i5[22:0]}),
              .i3({i2[1], i5[22:0], 1'b0}),
              .o1(o21[24:0]));
 m_18 inst_107(.i1(m121),
              .i2(i11[35:0]),
              .i3(i10[35:0]),
              .o1(m112[35:0]));
 m_8 inst_108(.i1(m121),
             .i2(m81),
             .i3(i5[31]),
             .o1(m123));
 m_8 inst_109(.i1(m121),
             .i2(m55),
             .i3(i5[31]),
             .o1(m76));
 m_16 inst_110(.i1(i3[1]),
              .i2(m106[31:0]),
              .i3({m112[26:23], m106[31:4]}),
              .o1(m85[31:0]));
 m_17 inst_111(.i1(i3[1]),
              .i2(10'b0010011110),
              .i3({1'b0, m112[35:27]}),
              .o1(o9[9:0]));
 m_5 inst_112(.i1(m28),
             .i2({m112[35:3], m29}),
             .i3({m112[35:27], m112[25:2], m30}),
             .o1(o4[33:0]));
 m_16 inst_113(.i1(o19),
              .i2({m85[15:0], 16'b0000000000000000}),
              .i3(m85[31:0]),
              .o1(m86[31:0]));
 m_15 inst_114(.i1(o18),
              .i2({m86[23:0], 8'b00000000}),
              .i3(m86[31:0]),
              .o1(o5[31:0]));
 m_16 inst_115(.i1(m120),
              .i2({i7[27:0], 4'b0000}),
              .i3(i7[31:0]),
              .o1(m87[31:0]));
 m_15 inst_116(.i1(m119),
              .i2({m87[29:0], 2'b00}),
              .i3(m87[31:0]),
              .o1(m88[31:0]));
 m_6 inst_117(.i1(m88[31]),
             .i2(m88[31:0]),
             .i3({m88[30:0], 1'b0}),
             .o1(m89[31:0]));
 m_14 inst_118(.i1(m18),
              .i2(i12[1:0]),
              .i3({m89[7], m31}),
              .o1(m102[1:0]));
 m_8 inst_119(.i1(i3[1]),
             .i2(m105[31]),
             .i3(m123),
             .o1(o10));
 m_13 inst_120(.i1(i14),
              .i2({i19, i16, 1'b0, i6[33:0]}),
              .i3({i19, i16, m99[9:0], m89[30:8], m102[1:0]}),
              .o1(m108[36:0]));
 m_10 inst_121(.i1(m32),
              .i2(5'b11111),
              .i3(m98[4:0]),
              .o1(m115[4:0]));
 m_10 inst_122(.i1(m33),
              .i2(5'b11111),
              .i3(m97[4:0]),
              .o1(m116[4:0]));
 m_12 inst_123(.i1(m98[8]),
              .i2({i4[30:23], 1'b1, i4[22:0]}),
              .i3({i5[30:23], 1'b1, i5[22:0]}),
              .o1(o17[31:0]));
 m_11 inst_124(.i1(m98[8]),
              .i2({i2[1], i5[22:0]}),
              .i3({i2[0], i4[22:0]}),
              .o1(m107[23:0]));
 m_11 inst_125(.i1(m100),
              .i2(24'b000000000000000000000000),
              .i3({i2[0], i4[22:0]}),
              .o1(m77[23:0]));
 m_11 inst_126(.i1(i3[1]),
              .i2(m77[23:0]),
              .i3(m107[23:0]),
              .o1(m111[23:0]));
 m_10 inst_127(.i1(m98[8]),
              .i2(m116[4:0]),
              .i3(m115[4:0]),
              .o1(m78[4:0]));
 m_10 inst_128(.i1(i3[1]),
              .i2(m113[4:0]),
              .i3(m78[4:0]),
              .o1(m117[4:0]));
 m_9 inst_129(.i1(m117[4]),
             .i2({16'b0000000000000000, m111[23:8], m34}),
             .i3({15'b000000000000000, m111[23:8], 2'b00}),
             .o1(m90[32:0]));
 m_9 inst_130(.i1(m117[3]),
             .i2({8'b00000000, m90[32:9], m35}),
             .i3(m90[32:0]),
             .o1(m91[32:0]));
 m_9 inst_131(.i1(m117[2]),
             .i2({4'b0000, m91[32:5], m36}),
             .i3(m91[32:0]),
             .o1(m92[32:0]));
 m_7 inst_132(.i1(m117[1]),
             .i2({2'b00, m92[32:3], m37}),
             .i3(m92[32:0]),
             .o1(m93[32:0]));
 m_9 inst_133(.i1(m117[0]),
             .i2({1'b0, m93[32:2], m38}),
             .i3(m93[32:0]),
             .o1({o14[27:2], m94[4:0], o14[1:0]}));
 m_8 inst_134(.i1(i4[31]),
             .i2(m11),
             .i3(1'b0),
             .o1(m79));
 m_7 inst_135(.i1(i4[31]),
             .i2({2'b11, m63[30:0]}),
             .i3({2'b00, o14[27:2], m94[4:0]}),
             .o1(m80[32:0]));
 m_6 inst_136(.i1(m104),
             .i2(32'b10000000000000000000000000000000),
             .i3(m101[31:0]),
             .o1(o3[31:0]));
 m_5 inst_137(.i1(m42),
             .i2({i18[35:3], m43}),
             .i3({i18[35:27], i18[25:2], m44}),
             .o1(m122[33:0]));
 m_5 inst_138(.i1(i18[26]),
             .i2({i18[35:27], i18[25:2], m45}),
             .i3({i18[35], m96[7:0], i18[24:0]}),
             .o1(m124[33:0]));
 m_4 inst_139(.i1(m59),
             .i2({m125, m123, 1'b0, m124[33:0]}),
             .i3({1'b0, m123, 1'b0, m122[33:0]}),
             .o1(o6[36:0]));
 m_3 inst_140(.i1(i17),
             .i2(m108[36:0]),
             .i3(i8[36:0]),
             .o1(o1[36:0]));
 m_2 inst_141(.i1(i3[0]),
             .i2(i4[31]),
             .o1(m81));
 m_2 inst_142(.i1(i4[31]),
             .i2(i5[31]),
             .o1(m82));
 m_2 inst_143(.i1(i3[0]),
             .i2(m82),
             .o1(m59));
 m_2 inst_144(.i1(i4[31]),
             .i2(m67),
             .o1(m83));
 m_1 inst_145(.i1({m105[31], m105[31], m105[31], m105[31], m105[31], m105[31], m105[31], m105[31], m105[31], m105[31], m105[31], m105[31], m105[31], m105[31], m105[31], m105[31], m105[31], m105[31], m105[31], m105[31], m105[31], m105[31], m105[31], m105[31], m105[31], m105[31], m105[31], m105[31], m105[31], m105[31], m105[31], m105[31]}),
             .i2(m105[31:0]),
             .o1(m84[31:0]));
 m inst_146(.i1(o15),
           .o1(m126));
 endmodule

 module m_53 (
    input [32 : 0] i1,
    input [32 : 0] i2,
    output [32 : 0] o1
 );
 assign o1 = i1[32:0] + i2[32:0];
 endmodule

 module m_52 (
    input [31 : 0] i1,
    input [31 : 0] i2,
    output [31 : 0] o1
 );
 assign o1 = i1[31:0] + i2[31:0];
 endmodule

 module m_51 (
    input i1,
    input i2,
    output o1
 );
 assign o1 = i1 & i2;
 endmodule

 module m_50 (
    input [31 : 0] i1,
    output o1
 );
 assign o1 = i1[31:0] == 32'b11001111000000000000000000000000;
 endmodule

 module m_49 (
    input [8 : 0] i1,
    output o1
 );
 assign o1 = i1[8:0] == 9'b111111111;
 endmodule

 module m_48 (
    input [31 : 0] i1,
    input [31 : 0] i2,
    output o1
 );
 assign o1 = i1[31:0] == i2[31:0];
 endmodule

 module m_47 (
    input [15 : 0] i1,
    output o1
 );
 assign o1 = i1[15:0] == 16'b0000000000000000;
 endmodule

 module m_46 (
    input [7 : 0] i1,
    output o1
 );
 assign o1 = i1[7:0] == 8'b00000000;
 endmodule

 module m_45 (
    input [3 : 0] i1,
    output o1
 );
 assign o1 = i1[3:0] == 4'b0000;
 endmodule

 module m_44 (
    input [31 : 0] i1,
    output o1
 );
 assign o1 = i1[31:0] == 32'b00000000000000000000000000000000;
 endmodule

 module m_43 (
    input [1 : 0] i1,
    output o1
 );
 assign o1 = i1[1:0] == 2'b10;
 endmodule

 module m_42 (
    input [2 : 0] i1,
    output o1
 );
 assign o1 = i1[2:0] == 3'b110;
 endmodule

 module m_41 (
    input [1 : 0] i1,
    output o1
 );
 assign o1 = i1[1:0] == 2'b11;
 endmodule

 module m_40 (
    input [26 : 0] i1,
    output o1
 );
 assign o1 = i1[26:0] == 27'b000000000000000000000000000;
 endmodule

 module m_39 (
    input [3 : 0] i1,
    output o1
 );
 assign o1 = ~(i1[3:0] == 4'b0000);
 endmodule

 module m_38 (
    input [7 : 0] i1,
    output o1
 );
 assign o1 = ~(i1[7:0] == 8'b00000000);
 endmodule

 module m_37 (
    input [8 : 0] i1,
    output o1
 );
 assign o1 = ~(i1[8:0] == 9'b000000000);
 endmodule

 module m_36 (
    input [4 : 0] i1,
    output o1
 );
 assign o1 = ~(i1[4:0] == 5'b00000);
 endmodule

 module m_35 (
    input [6 : 0] i1,
    output o1
 );
 assign o1 = ~(i1[6:0] == 7'b0000000);
 endmodule

 module m_34 (
    input i1,
    input i2,
    output o1
 );
 assign o1 = ~(i1 == i2);
 endmodule

 module m_33 (
    input [2 : 0] i1,
    output o1
 );
 assign o1 = ~(i1[2:0] == 3'b000);
 endmodule

 module m_32 (
    input [1 : 0] i1,
    output o1
 );
 assign o1 = ~(i1[1:0] == 2'b00);
 endmodule

 module m_31 (
    input i1,
    output o1
 );
 assign o1 = ~(i1);
 endmodule

 module m_30 (
    input [30 : 0] i1,
    output [30 : 0] o1
 );
 assign o1 = ~(i1[30:0]);
 endmodule

 module m_29 (
    input [9 : 0] i1,
    input [9 : 0] i2,
    output [9 : 0] o1
 );
 assign o1 = i1[9:0] | i2[9:0];
 endmodule

 module m_28 (
    input i1,
    input i2,
    output o1
 );
 assign o1 = i1 | i2;
 endmodule

 module m_27 (
    input i1,
    input i2,
    input i3,
    input i4,
    input i5,
    output o1
 );
 assign o1 = i1 ? i2 : i3 ? i4 : i5;
 endmodule

 module m_26 (
    input i1,
    input [31 : 0] i2,
    input i3,
    input [31 : 0] i4,
    input [31 : 0] i5,
    output [31 : 0] o1
 );
 assign o1 = i1 ? i2[31:0] : i3 ? i4[31:0] : i5[31:0];
 endmodule

 module m_25 (
    input [1 : 0] i1,
    output o1
 );
 assign o1 = i1[1:0] == 2'b01;
 endmodule

 module m_24 (
    input [1 : 0] i1,
    output o1
 );
 assign o1 = i1[1:0] == 2'b00;
 endmodule

 module m_23 (
    input [23 : 0] i1,
    input [23 : 0] i2,
    output [23 : 0] o1
 );
 assign o1 = i1[23:0] - i2[23:0];
 endmodule

 module m_22 (
    input [9 : 0] i1,
    input [9 : 0] i2,
    output [9 : 0] o1
 );
 assign o1 = i1[9:0] - i2[9:0];
 endmodule

 module m_21 (
    input [8 : 0] i1,
    input [8 : 0] i2,
    output [8 : 0] o1
 );
 assign o1 = i1[8:0] - i2[8:0];
 endmodule

 module m_20 (
    input [7 : 0] i1,
    input [7 : 0] i2,
    output [7 : 0] o1
 );
 assign o1 = i1[7:0] - i2[7:0];
 endmodule

 module m_19 (
    input i1,
    input [24 : 0] i2,
    input [24 : 0] i3,
    output [24 : 0] o1
 );
 assign o1 = i1 ? i2[24:0] : i3[24:0];
 endmodule

 module m_18 (
    input i1,
    input [35 : 0] i2,
    input [35 : 0] i3,
    output [35 : 0] o1
 );
 assign o1 = i1 ? i2[35:0] : i3[35:0];
 endmodule

 module m_17 (
    input i1,
    input [9 : 0] i2,
    input [9 : 0] i3,
    output [9 : 0] o1
 );
 assign o1 = i1 ? i2[9:0] : i3[9:0];
 endmodule

 module m_16 (
    input i1,
    input [31 : 0] i2,
    input [31 : 0] i3,
    output [31 : 0] o1
 );
 assign o1 = i1 ? i2[31:0] : i3[31:0];
 endmodule

 module m_15 (
    input i1,
    input [31 : 0] i2,
    input [31 : 0] i3,
    output [31 : 0] o1
 );
 assign o1 = i1 ? i2[31:0] : i3[31:0];
 endmodule

 module m_14 (
    input i1,
    input [1 : 0] i2,
    input [1 : 0] i3,
    output [1 : 0] o1
 );
 assign o1 = i1 ? i2[1:0] : i3[1:0];
 endmodule

 module m_13 (
    input i1,
    input [36 : 0] i2,
    input [36 : 0] i3,
    output [36 : 0] o1
 );
 assign o1 = i1 ? i2[36:0] : i3[36:0];
 endmodule

 module m_12 (
    input i1,
    input [31 : 0] i2,
    input [31 : 0] i3,
    output [31 : 0] o1
 );
 assign o1 = i1 ? i2[31:0] : i3[31:0];
 endmodule

 module m_11 (
    input i1,
    input [23 : 0] i2,
    input [23 : 0] i3,
    output [23 : 0] o1
 );
 assign o1 = i1 ? i2[23:0] : i3[23:0];
 endmodule

 module m_10 (
    input i1,
    input [4 : 0] i2,
    input [4 : 0] i3,
    output [4 : 0] o1
 );
 assign o1 = i1 ? i2[4:0] : i3[4:0];
 endmodule

 module m_9 (
    input i1,
    input [32 : 0] i2,
    input [32 : 0] i3,
    output [32 : 0] o1
 );
 assign o1 = i1 ? i2[32:0] : i3[32:0];
 endmodule

 module m_8 (
    input i1,
    input i2,
    input i3,
    output o1
 );
 assign o1 = i1 ? i2 : i3;
 endmodule

 module m_7 (
    input i1,
    input [32 : 0] i2,
    input [32 : 0] i3,
    output [32 : 0] o1
 );
 assign o1 = i1 ? i2[32:0] : i3[32:0];
 endmodule

 module m_6 (
    input i1,
    input [31 : 0] i2,
    input [31 : 0] i3,
    output [31 : 0] o1
 );
 assign o1 = i1 ? i2[31:0] : i3[31:0];
 endmodule

 module m_5 (
    input i1,
    input [33 : 0] i2,
    input [33 : 0] i3,
    output [33 : 0] o1
 );
 assign o1 = i1 ? i2[33:0] : i3[33:0];
 endmodule

 module m_4 (
    input i1,
    input [36 : 0] i2,
    input [36 : 0] i3,
    output [36 : 0] o1
 );
 assign o1 = i1 ? i2[36:0] : i3[36:0];
 endmodule

 module m_3 (
    input i1,
    input [36 : 0] i2,
    input [36 : 0] i3,
    output [36 : 0] o1
 );
 assign o1 = i1 ? i2[36:0] : i3[36:0];
 endmodule

 module m_2 (
    input i1,
    input i2,
    output o1
 );
 assign o1 = ~(i1) & i2 | i1 & ~(i2);
 endmodule

 module m_1 (
    input [31 : 0] i1,
    input [31 : 0] i2,
    output [31 : 0] o1
 );
 assign o1 = ~(i1[31:0]) & i2[31:0] | i1[31:0] & ~(i2[31:0]);
 endmodule

 module m (
    input i1,
    output o1
 );
 assign o1 = i1;
 endmodule

